library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.types.all;

package prog_mem is

	constant PROG_SIZE : integer := 96956;

	constant PROG_DATA : mem_type(0 to PROG_SIZE/4-1) := (
		16#0000# => X"93000000",
		16#0001# => X"13010000",
		16#0002# => X"93010000",
		16#0003# => X"13020000",
		16#0004# => X"93020000",
		16#0005# => X"13030000",
		16#0006# => X"93030000",
		16#0007# => X"13040000",
		16#0008# => X"93040000",
		16#0009# => X"13050000",
		16#000a# => X"93050000",
		16#000b# => X"13060000",
		16#000c# => X"93060000",
		16#000d# => X"13070000",
		16#000e# => X"93070000",
		16#000f# => X"13080000",
		16#0010# => X"93080000",
		16#0011# => X"13090000",
		16#0012# => X"93090000",
		16#0013# => X"130a0000",
		16#0014# => X"930a0000",
		16#0015# => X"130b0000",
		16#0016# => X"930b0000",
		16#0017# => X"130c0000",
		16#0018# => X"930c0000",
		16#0019# => X"130d0000",
		16#001a# => X"930d0000",
		16#001b# => X"130e0000",
		16#001c# => X"930e0000",
		16#001d# => X"130f0000",
		16#001e# => X"930f0000",
		16#001f# => X"732540f1",
		16#0020# => X"63180502",
		16#0021# => X"73a00230",
		16#0022# => X"93021000",
		16#0023# => X"9392f201",
		16#0024# => X"63ca0200",
		16#0025# => X"13051000",
		16#0026# => X"97120000",
		16#0027# => X"23a4a2f6",
		16#0028# => X"6ff05fff",
		16#0029# => X"97020000",
		16#002a# => X"9382c203",
		16#002b# => X"73905230",
		16#002c# => X"97610100",
		16#002d# => X"93818196",
		16#002e# => X"17820100",
		16#002f# => X"130272f8",
		16#0030# => X"1302c203",
		16#0031# => X"137202fc",
		16#0032# => X"13161501",
		16#0033# => X"3302c200",
		16#0034# => X"13011500",
		16#0035# => X"13111101",
		16#0036# => X"33014100",
		16#0037# => X"6fd00001",
		16#0038# => X"130101ef",
		16#0039# => X"23221100",
		16#003a# => X"23242100",
		16#003b# => X"23263100",
		16#003c# => X"23284100",
		16#003d# => X"232a5100",
		16#003e# => X"232c6100",
		16#003f# => X"232e7100",
		16#0040# => X"23208102",
		16#0041# => X"23229102",
		16#0042# => X"2324a102",
		16#0043# => X"2326b102",
		16#0044# => X"2328c102",
		16#0045# => X"232ad102",
		16#0046# => X"232ce102",
		16#0047# => X"232ef102",
		16#0048# => X"23200105",
		16#0049# => X"23221105",
		16#004a# => X"23242105",
		16#004b# => X"23263105",
		16#004c# => X"23284105",
		16#004d# => X"232a5105",
		16#004e# => X"232c6105",
		16#004f# => X"232e7105",
		16#0050# => X"23208107",
		16#0051# => X"23229107",
		16#0052# => X"2324a107",
		16#0053# => X"2326b107",
		16#0054# => X"2328c107",
		16#0055# => X"232ad107",
		16#0056# => X"232ce107",
		16#0057# => X"232ef107",
		16#0058# => X"73252034",
		16#0059# => X"f3251034",
		16#005a# => X"13060100",
		16#005b# => X"73101534",
		16#005c# => X"83204100",
		16#005d# => X"03218100",
		16#005e# => X"8321c100",
		16#005f# => X"03220101",
		16#0060# => X"83224101",
		16#0061# => X"03238101",
		16#0062# => X"8323c101",
		16#0063# => X"03240102",
		16#0064# => X"83244102",
		16#0065# => X"03258102",
		16#0066# => X"8325c102",
		16#0067# => X"03260103",
		16#0068# => X"83264103",
		16#0069# => X"03278103",
		16#006a# => X"8327c103",
		16#006b# => X"03280104",
		16#006c# => X"83284104",
		16#006d# => X"03298104",
		16#006e# => X"8329c104",
		16#006f# => X"032a0105",
		16#0070# => X"832a4105",
		16#0071# => X"032b8105",
		16#0072# => X"832bc105",
		16#0073# => X"032c0106",
		16#0074# => X"832c4106",
		16#0075# => X"032d8106",
		16#0076# => X"832dc106",
		16#0077# => X"032e0107",
		16#0078# => X"832e4107",
		16#0079# => X"032f8107",
		16#007a# => X"832fc107",
		16#007b# => X"13010111",
		16#007c# => X"67800000",
		16#007d# => X"00000000",
		16#007e# => X"00000000",
		16#007f# => X"00000000",
		16#0080# => X"00000000",
		16#0081# => X"00000000",
		16#0082# => X"00000000",
		16#0083# => X"00000000",
		16#0084# => X"00000000",
		16#0085# => X"00000000",
		16#0086# => X"00000000",
		16#0087# => X"00000000",
		16#0088# => X"00000000",
		16#0089# => X"00000000",
		16#008a# => X"00000000",
		16#008b# => X"00000000",
		16#008c# => X"00000000",
		16#008d# => X"00000000",
		16#008e# => X"00000000",
		16#008f# => X"00000000",
		16#0090# => X"00000000",
		16#0091# => X"00000000",
		16#0092# => X"00000000",
		16#0093# => X"00000000",
		16#0094# => X"00000000",
		16#0095# => X"00000000",
		16#0096# => X"00000000",
		16#0097# => X"00000000",
		16#0098# => X"00000000",
		16#0099# => X"00000000",
		16#009a# => X"00000000",
		16#009b# => X"00000000",
		16#009c# => X"00000000",
		16#009d# => X"00000000",
		16#009e# => X"00000000",
		16#009f# => X"00000000",
		16#00a0# => X"00000000",
		16#00a1# => X"00000000",
		16#00a2# => X"00000000",
		16#00a3# => X"00000000",
		16#00a4# => X"00000000",
		16#00a5# => X"00000000",
		16#00a6# => X"00000000",
		16#00a7# => X"00000000",
		16#00a8# => X"00000000",
		16#00a9# => X"00000000",
		16#00aa# => X"00000000",
		16#00ab# => X"00000000",
		16#00ac# => X"00000000",
		16#00ad# => X"00000000",
		16#00ae# => X"00000000",
		16#00af# => X"00000000",
		16#00b0# => X"00000000",
		16#00b1# => X"00000000",
		16#00b2# => X"00000000",
		16#00b3# => X"00000000",
		16#00b4# => X"00000000",
		16#00b5# => X"00000000",
		16#00b6# => X"00000000",
		16#00b7# => X"00000000",
		16#00b8# => X"00000000",
		16#00b9# => X"00000000",
		16#00ba# => X"00000000",
		16#00bb# => X"00000000",
		16#00bc# => X"00000000",
		16#00bd# => X"00000000",
		16#00be# => X"00000000",
		16#00bf# => X"00000000",
		16#00c0# => X"00000000",
		16#00c1# => X"00000000",
		16#00c2# => X"00000000",
		16#00c3# => X"00000000",
		16#00c4# => X"00000000",
		16#00c5# => X"00000000",
		16#00c6# => X"00000000",
		16#00c7# => X"00000000",
		16#00c8# => X"00000000",
		16#00c9# => X"00000000",
		16#00ca# => X"00000000",
		16#00cb# => X"00000000",
		16#00cc# => X"00000000",
		16#00cd# => X"00000000",
		16#00ce# => X"00000000",
		16#00cf# => X"00000000",
		16#00d0# => X"00000000",
		16#00d1# => X"00000000",
		16#00d2# => X"00000000",
		16#00d3# => X"00000000",
		16#00d4# => X"00000000",
		16#00d5# => X"00000000",
		16#00d6# => X"00000000",
		16#00d7# => X"00000000",
		16#00d8# => X"00000000",
		16#00d9# => X"00000000",
		16#00da# => X"00000000",
		16#00db# => X"00000000",
		16#00dc# => X"00000000",
		16#00dd# => X"00000000",
		16#00de# => X"00000000",
		16#00df# => X"00000000",
		16#00e0# => X"00000000",
		16#00e1# => X"00000000",
		16#00e2# => X"00000000",
		16#00e3# => X"00000000",
		16#00e4# => X"00000000",
		16#00e5# => X"00000000",
		16#00e6# => X"00000000",
		16#00e7# => X"00000000",
		16#00e8# => X"00000000",
		16#00e9# => X"00000000",
		16#00ea# => X"00000000",
		16#00eb# => X"00000000",
		16#00ec# => X"00000000",
		16#00ed# => X"00000000",
		16#00ee# => X"00000000",
		16#00ef# => X"00000000",
		16#00f0# => X"00000000",
		16#00f1# => X"00000000",
		16#00f2# => X"00000000",
		16#00f3# => X"00000000",
		16#00f4# => X"00000000",
		16#00f5# => X"00000000",
		16#00f6# => X"00000000",
		16#00f7# => X"00000000",
		16#00f8# => X"00000000",
		16#00f9# => X"00000000",
		16#00fa# => X"00000000",
		16#00fb# => X"00000000",
		16#00fc# => X"00000000",
		16#00fd# => X"00000000",
		16#00fe# => X"00000000",
		16#00ff# => X"00000000",
		16#0100# => X"00000000",
		16#0101# => X"00000000",
		16#0102# => X"00000000",
		16#0103# => X"00000000",
		16#0104# => X"00000000",
		16#0105# => X"00000000",
		16#0106# => X"00000000",
		16#0107# => X"00000000",
		16#0108# => X"00000000",
		16#0109# => X"00000000",
		16#010a# => X"00000000",
		16#010b# => X"00000000",
		16#010c# => X"00000000",
		16#010d# => X"00000000",
		16#010e# => X"00000000",
		16#010f# => X"00000000",
		16#0110# => X"00000000",
		16#0111# => X"00000000",
		16#0112# => X"00000000",
		16#0113# => X"00000000",
		16#0114# => X"00000000",
		16#0115# => X"00000000",
		16#0116# => X"00000000",
		16#0117# => X"00000000",
		16#0118# => X"00000000",
		16#0119# => X"00000000",
		16#011a# => X"00000000",
		16#011b# => X"00000000",
		16#011c# => X"00000000",
		16#011d# => X"00000000",
		16#011e# => X"00000000",
		16#011f# => X"00000000",
		16#0120# => X"00000000",
		16#0121# => X"00000000",
		16#0122# => X"00000000",
		16#0123# => X"00000000",
		16#0124# => X"00000000",
		16#0125# => X"00000000",
		16#0126# => X"00000000",
		16#0127# => X"00000000",
		16#0128# => X"00000000",
		16#0129# => X"00000000",
		16#012a# => X"00000000",
		16#012b# => X"00000000",
		16#012c# => X"00000000",
		16#012d# => X"00000000",
		16#012e# => X"00000000",
		16#012f# => X"00000000",
		16#0130# => X"00000000",
		16#0131# => X"00000000",
		16#0132# => X"00000000",
		16#0133# => X"00000000",
		16#0134# => X"00000000",
		16#0135# => X"00000000",
		16#0136# => X"00000000",
		16#0137# => X"00000000",
		16#0138# => X"00000000",
		16#0139# => X"00000000",
		16#013a# => X"00000000",
		16#013b# => X"00000000",
		16#013c# => X"00000000",
		16#013d# => X"00000000",
		16#013e# => X"00000000",
		16#013f# => X"00000000",
		16#0140# => X"00000000",
		16#0141# => X"00000000",
		16#0142# => X"00000000",
		16#0143# => X"00000000",
		16#0144# => X"00000000",
		16#0145# => X"00000000",
		16#0146# => X"00000000",
		16#0147# => X"00000000",
		16#0148# => X"00000000",
		16#0149# => X"00000000",
		16#014a# => X"00000000",
		16#014b# => X"00000000",
		16#014c# => X"00000000",
		16#014d# => X"00000000",
		16#014e# => X"00000000",
		16#014f# => X"00000000",
		16#0150# => X"00000000",
		16#0151# => X"00000000",
		16#0152# => X"00000000",
		16#0153# => X"00000000",
		16#0154# => X"00000000",
		16#0155# => X"00000000",
		16#0156# => X"00000000",
		16#0157# => X"00000000",
		16#0158# => X"00000000",
		16#0159# => X"00000000",
		16#015a# => X"00000000",
		16#015b# => X"00000000",
		16#015c# => X"00000000",
		16#015d# => X"00000000",
		16#015e# => X"00000000",
		16#015f# => X"00000000",
		16#0160# => X"00000000",
		16#0161# => X"00000000",
		16#0162# => X"00000000",
		16#0163# => X"00000000",
		16#0164# => X"00000000",
		16#0165# => X"00000000",
		16#0166# => X"00000000",
		16#0167# => X"00000000",
		16#0168# => X"00000000",
		16#0169# => X"00000000",
		16#016a# => X"00000000",
		16#016b# => X"00000000",
		16#016c# => X"00000000",
		16#016d# => X"00000000",
		16#016e# => X"00000000",
		16#016f# => X"00000000",
		16#0170# => X"00000000",
		16#0171# => X"00000000",
		16#0172# => X"00000000",
		16#0173# => X"00000000",
		16#0174# => X"00000000",
		16#0175# => X"00000000",
		16#0176# => X"00000000",
		16#0177# => X"00000000",
		16#0178# => X"00000000",
		16#0179# => X"00000000",
		16#017a# => X"00000000",
		16#017b# => X"00000000",
		16#017c# => X"00000000",
		16#017d# => X"00000000",
		16#017e# => X"00000000",
		16#017f# => X"00000000",
		16#0180# => X"00000000",
		16#0181# => X"00000000",
		16#0182# => X"00000000",
		16#0183# => X"00000000",
		16#0184# => X"00000000",
		16#0185# => X"00000000",
		16#0186# => X"00000000",
		16#0187# => X"00000000",
		16#0188# => X"00000000",
		16#0189# => X"00000000",
		16#018a# => X"00000000",
		16#018b# => X"00000000",
		16#018c# => X"00000000",
		16#018d# => X"00000000",
		16#018e# => X"00000000",
		16#018f# => X"00000000",
		16#0190# => X"00000000",
		16#0191# => X"00000000",
		16#0192# => X"00000000",
		16#0193# => X"00000000",
		16#0194# => X"00000000",
		16#0195# => X"00000000",
		16#0196# => X"00000000",
		16#0197# => X"00000000",
		16#0198# => X"00000000",
		16#0199# => X"00000000",
		16#019a# => X"00000000",
		16#019b# => X"00000000",
		16#019c# => X"00000000",
		16#019d# => X"00000000",
		16#019e# => X"00000000",
		16#019f# => X"00000000",
		16#01a0# => X"00000000",
		16#01a1# => X"00000000",
		16#01a2# => X"00000000",
		16#01a3# => X"00000000",
		16#01a4# => X"00000000",
		16#01a5# => X"00000000",
		16#01a6# => X"00000000",
		16#01a7# => X"00000000",
		16#01a8# => X"00000000",
		16#01a9# => X"00000000",
		16#01aa# => X"00000000",
		16#01ab# => X"00000000",
		16#01ac# => X"00000000",
		16#01ad# => X"00000000",
		16#01ae# => X"00000000",
		16#01af# => X"00000000",
		16#01b0# => X"00000000",
		16#01b1# => X"00000000",
		16#01b2# => X"00000000",
		16#01b3# => X"00000000",
		16#01b4# => X"00000000",
		16#01b5# => X"00000000",
		16#01b6# => X"00000000",
		16#01b7# => X"00000000",
		16#01b8# => X"00000000",
		16#01b9# => X"00000000",
		16#01ba# => X"00000000",
		16#01bb# => X"00000000",
		16#01bc# => X"00000000",
		16#01bd# => X"00000000",
		16#01be# => X"00000000",
		16#01bf# => X"00000000",
		16#01c0# => X"00000000",
		16#01c1# => X"00000000",
		16#01c2# => X"00000000",
		16#01c3# => X"00000000",
		16#01c4# => X"00000000",
		16#01c5# => X"00000000",
		16#01c6# => X"00000000",
		16#01c7# => X"00000000",
		16#01c8# => X"00000000",
		16#01c9# => X"00000000",
		16#01ca# => X"00000000",
		16#01cb# => X"00000000",
		16#01cc# => X"00000000",
		16#01cd# => X"00000000",
		16#01ce# => X"00000000",
		16#01cf# => X"00000000",
		16#01d0# => X"00000000",
		16#01d1# => X"00000000",
		16#01d2# => X"00000000",
		16#01d3# => X"00000000",
		16#01d4# => X"00000000",
		16#01d5# => X"00000000",
		16#01d6# => X"00000000",
		16#01d7# => X"00000000",
		16#01d8# => X"00000000",
		16#01d9# => X"00000000",
		16#01da# => X"00000000",
		16#01db# => X"00000000",
		16#01dc# => X"00000000",
		16#01dd# => X"00000000",
		16#01de# => X"00000000",
		16#01df# => X"00000000",
		16#01e0# => X"00000000",
		16#01e1# => X"00000000",
		16#01e2# => X"00000000",
		16#01e3# => X"00000000",
		16#01e4# => X"00000000",
		16#01e5# => X"00000000",
		16#01e6# => X"00000000",
		16#01e7# => X"00000000",
		16#01e8# => X"00000000",
		16#01e9# => X"00000000",
		16#01ea# => X"00000000",
		16#01eb# => X"00000000",
		16#01ec# => X"00000000",
		16#01ed# => X"00000000",
		16#01ee# => X"00000000",
		16#01ef# => X"00000000",
		16#01f0# => X"00000000",
		16#01f1# => X"00000000",
		16#01f2# => X"00000000",
		16#01f3# => X"00000000",
		16#01f4# => X"00000000",
		16#01f5# => X"00000000",
		16#01f6# => X"00000000",
		16#01f7# => X"00000000",
		16#01f8# => X"00000000",
		16#01f9# => X"00000000",
		16#01fa# => X"00000000",
		16#01fb# => X"00000000",
		16#01fc# => X"00000000",
		16#01fd# => X"00000000",
		16#01fe# => X"00000000",
		16#01ff# => X"00000000",
		16#0200# => X"00000000",
		16#0201# => X"00000000",
		16#0202# => X"00000000",
		16#0203# => X"00000000",
		16#0204# => X"00000000",
		16#0205# => X"00000000",
		16#0206# => X"00000000",
		16#0207# => X"00000000",
		16#0208# => X"00000000",
		16#0209# => X"00000000",
		16#020a# => X"00000000",
		16#020b# => X"00000000",
		16#020c# => X"00000000",
		16#020d# => X"00000000",
		16#020e# => X"00000000",
		16#020f# => X"00000000",
		16#0210# => X"00000000",
		16#0211# => X"00000000",
		16#0212# => X"00000000",
		16#0213# => X"00000000",
		16#0214# => X"00000000",
		16#0215# => X"00000000",
		16#0216# => X"00000000",
		16#0217# => X"00000000",
		16#0218# => X"00000000",
		16#0219# => X"00000000",
		16#021a# => X"00000000",
		16#021b# => X"00000000",
		16#021c# => X"00000000",
		16#021d# => X"00000000",
		16#021e# => X"00000000",
		16#021f# => X"00000000",
		16#0220# => X"00000000",
		16#0221# => X"00000000",
		16#0222# => X"00000000",
		16#0223# => X"00000000",
		16#0224# => X"00000000",
		16#0225# => X"00000000",
		16#0226# => X"00000000",
		16#0227# => X"00000000",
		16#0228# => X"00000000",
		16#0229# => X"00000000",
		16#022a# => X"00000000",
		16#022b# => X"00000000",
		16#022c# => X"00000000",
		16#022d# => X"00000000",
		16#022e# => X"00000000",
		16#022f# => X"00000000",
		16#0230# => X"00000000",
		16#0231# => X"00000000",
		16#0232# => X"00000000",
		16#0233# => X"00000000",
		16#0234# => X"00000000",
		16#0235# => X"00000000",
		16#0236# => X"00000000",
		16#0237# => X"00000000",
		16#0238# => X"00000000",
		16#0239# => X"00000000",
		16#023a# => X"00000000",
		16#023b# => X"00000000",
		16#023c# => X"00000000",
		16#023d# => X"00000000",
		16#023e# => X"00000000",
		16#023f# => X"00000000",
		16#0240# => X"00000000",
		16#0241# => X"00000000",
		16#0242# => X"00000000",
		16#0243# => X"00000000",
		16#0244# => X"00000000",
		16#0245# => X"00000000",
		16#0246# => X"00000000",
		16#0247# => X"00000000",
		16#0248# => X"00000000",
		16#0249# => X"00000000",
		16#024a# => X"00000000",
		16#024b# => X"00000000",
		16#024c# => X"00000000",
		16#024d# => X"00000000",
		16#024e# => X"00000000",
		16#024f# => X"00000000",
		16#0250# => X"00000000",
		16#0251# => X"00000000",
		16#0252# => X"00000000",
		16#0253# => X"00000000",
		16#0254# => X"00000000",
		16#0255# => X"00000000",
		16#0256# => X"00000000",
		16#0257# => X"00000000",
		16#0258# => X"00000000",
		16#0259# => X"00000000",
		16#025a# => X"00000000",
		16#025b# => X"00000000",
		16#025c# => X"00000000",
		16#025d# => X"00000000",
		16#025e# => X"00000000",
		16#025f# => X"00000000",
		16#0260# => X"00000000",
		16#0261# => X"00000000",
		16#0262# => X"00000000",
		16#0263# => X"00000000",
		16#0264# => X"00000000",
		16#0265# => X"00000000",
		16#0266# => X"00000000",
		16#0267# => X"00000000",
		16#0268# => X"00000000",
		16#0269# => X"00000000",
		16#026a# => X"00000000",
		16#026b# => X"00000000",
		16#026c# => X"00000000",
		16#026d# => X"00000000",
		16#026e# => X"00000000",
		16#026f# => X"00000000",
		16#0270# => X"00000000",
		16#0271# => X"00000000",
		16#0272# => X"00000000",
		16#0273# => X"00000000",
		16#0274# => X"00000000",
		16#0275# => X"00000000",
		16#0276# => X"00000000",
		16#0277# => X"00000000",
		16#0278# => X"00000000",
		16#0279# => X"00000000",
		16#027a# => X"00000000",
		16#027b# => X"00000000",
		16#027c# => X"00000000",
		16#027d# => X"00000000",
		16#027e# => X"00000000",
		16#027f# => X"00000000",
		16#0280# => X"00000000",
		16#0281# => X"00000000",
		16#0282# => X"00000000",
		16#0283# => X"00000000",
		16#0284# => X"00000000",
		16#0285# => X"00000000",
		16#0286# => X"00000000",
		16#0287# => X"00000000",
		16#0288# => X"00000000",
		16#0289# => X"00000000",
		16#028a# => X"00000000",
		16#028b# => X"00000000",
		16#028c# => X"00000000",
		16#028d# => X"00000000",
		16#028e# => X"00000000",
		16#028f# => X"00000000",
		16#0290# => X"00000000",
		16#0291# => X"00000000",
		16#0292# => X"00000000",
		16#0293# => X"00000000",
		16#0294# => X"00000000",
		16#0295# => X"00000000",
		16#0296# => X"00000000",
		16#0297# => X"00000000",
		16#0298# => X"00000000",
		16#0299# => X"00000000",
		16#029a# => X"00000000",
		16#029b# => X"00000000",
		16#029c# => X"00000000",
		16#029d# => X"00000000",
		16#029e# => X"00000000",
		16#029f# => X"00000000",
		16#02a0# => X"00000000",
		16#02a1# => X"00000000",
		16#02a2# => X"00000000",
		16#02a3# => X"00000000",
		16#02a4# => X"00000000",
		16#02a5# => X"00000000",
		16#02a6# => X"00000000",
		16#02a7# => X"00000000",
		16#02a8# => X"00000000",
		16#02a9# => X"00000000",
		16#02aa# => X"00000000",
		16#02ab# => X"00000000",
		16#02ac# => X"00000000",
		16#02ad# => X"00000000",
		16#02ae# => X"00000000",
		16#02af# => X"00000000",
		16#02b0# => X"00000000",
		16#02b1# => X"00000000",
		16#02b2# => X"00000000",
		16#02b3# => X"00000000",
		16#02b4# => X"00000000",
		16#02b5# => X"00000000",
		16#02b6# => X"00000000",
		16#02b7# => X"00000000",
		16#02b8# => X"00000000",
		16#02b9# => X"00000000",
		16#02ba# => X"00000000",
		16#02bb# => X"00000000",
		16#02bc# => X"00000000",
		16#02bd# => X"00000000",
		16#02be# => X"00000000",
		16#02bf# => X"00000000",
		16#02c0# => X"00000000",
		16#02c1# => X"00000000",
		16#02c2# => X"00000000",
		16#02c3# => X"00000000",
		16#02c4# => X"00000000",
		16#02c5# => X"00000000",
		16#02c6# => X"00000000",
		16#02c7# => X"00000000",
		16#02c8# => X"00000000",
		16#02c9# => X"00000000",
		16#02ca# => X"00000000",
		16#02cb# => X"00000000",
		16#02cc# => X"00000000",
		16#02cd# => X"00000000",
		16#02ce# => X"00000000",
		16#02cf# => X"00000000",
		16#02d0# => X"00000000",
		16#02d1# => X"00000000",
		16#02d2# => X"00000000",
		16#02d3# => X"00000000",
		16#02d4# => X"00000000",
		16#02d5# => X"00000000",
		16#02d6# => X"00000000",
		16#02d7# => X"00000000",
		16#02d8# => X"00000000",
		16#02d9# => X"00000000",
		16#02da# => X"00000000",
		16#02db# => X"00000000",
		16#02dc# => X"00000000",
		16#02dd# => X"00000000",
		16#02de# => X"00000000",
		16#02df# => X"00000000",
		16#02e0# => X"00000000",
		16#02e1# => X"00000000",
		16#02e2# => X"00000000",
		16#02e3# => X"00000000",
		16#02e4# => X"00000000",
		16#02e5# => X"00000000",
		16#02e6# => X"00000000",
		16#02e7# => X"00000000",
		16#02e8# => X"00000000",
		16#02e9# => X"00000000",
		16#02ea# => X"00000000",
		16#02eb# => X"00000000",
		16#02ec# => X"00000000",
		16#02ed# => X"00000000",
		16#02ee# => X"00000000",
		16#02ef# => X"00000000",
		16#02f0# => X"00000000",
		16#02f1# => X"00000000",
		16#02f2# => X"00000000",
		16#02f3# => X"00000000",
		16#02f4# => X"00000000",
		16#02f5# => X"00000000",
		16#02f6# => X"00000000",
		16#02f7# => X"00000000",
		16#02f8# => X"00000000",
		16#02f9# => X"00000000",
		16#02fa# => X"00000000",
		16#02fb# => X"00000000",
		16#02fc# => X"00000000",
		16#02fd# => X"00000000",
		16#02fe# => X"00000000",
		16#02ff# => X"00000000",
		16#0300# => X"00000000",
		16#0301# => X"00000000",
		16#0302# => X"00000000",
		16#0303# => X"00000000",
		16#0304# => X"00000000",
		16#0305# => X"00000000",
		16#0306# => X"00000000",
		16#0307# => X"00000000",
		16#0308# => X"00000000",
		16#0309# => X"00000000",
		16#030a# => X"00000000",
		16#030b# => X"00000000",
		16#030c# => X"00000000",
		16#030d# => X"00000000",
		16#030e# => X"00000000",
		16#030f# => X"00000000",
		16#0310# => X"00000000",
		16#0311# => X"00000000",
		16#0312# => X"00000000",
		16#0313# => X"00000000",
		16#0314# => X"00000000",
		16#0315# => X"00000000",
		16#0316# => X"00000000",
		16#0317# => X"00000000",
		16#0318# => X"00000000",
		16#0319# => X"00000000",
		16#031a# => X"00000000",
		16#031b# => X"00000000",
		16#031c# => X"00000000",
		16#031d# => X"00000000",
		16#031e# => X"00000000",
		16#031f# => X"00000000",
		16#0320# => X"00000000",
		16#0321# => X"00000000",
		16#0322# => X"00000000",
		16#0323# => X"00000000",
		16#0324# => X"00000000",
		16#0325# => X"00000000",
		16#0326# => X"00000000",
		16#0327# => X"00000000",
		16#0328# => X"00000000",
		16#0329# => X"00000000",
		16#032a# => X"00000000",
		16#032b# => X"00000000",
		16#032c# => X"00000000",
		16#032d# => X"00000000",
		16#032e# => X"00000000",
		16#032f# => X"00000000",
		16#0330# => X"00000000",
		16#0331# => X"00000000",
		16#0332# => X"00000000",
		16#0333# => X"00000000",
		16#0334# => X"00000000",
		16#0335# => X"00000000",
		16#0336# => X"00000000",
		16#0337# => X"00000000",
		16#0338# => X"00000000",
		16#0339# => X"00000000",
		16#033a# => X"00000000",
		16#033b# => X"00000000",
		16#033c# => X"00000000",
		16#033d# => X"00000000",
		16#033e# => X"00000000",
		16#033f# => X"00000000",
		16#0340# => X"00000000",
		16#0341# => X"00000000",
		16#0342# => X"00000000",
		16#0343# => X"00000000",
		16#0344# => X"00000000",
		16#0345# => X"00000000",
		16#0346# => X"00000000",
		16#0347# => X"00000000",
		16#0348# => X"00000000",
		16#0349# => X"00000000",
		16#034a# => X"00000000",
		16#034b# => X"00000000",
		16#034c# => X"00000000",
		16#034d# => X"00000000",
		16#034e# => X"00000000",
		16#034f# => X"00000000",
		16#0350# => X"00000000",
		16#0351# => X"00000000",
		16#0352# => X"00000000",
		16#0353# => X"00000000",
		16#0354# => X"00000000",
		16#0355# => X"00000000",
		16#0356# => X"00000000",
		16#0357# => X"00000000",
		16#0358# => X"00000000",
		16#0359# => X"00000000",
		16#035a# => X"00000000",
		16#035b# => X"00000000",
		16#035c# => X"00000000",
		16#035d# => X"00000000",
		16#035e# => X"00000000",
		16#035f# => X"00000000",
		16#0360# => X"00000000",
		16#0361# => X"00000000",
		16#0362# => X"00000000",
		16#0363# => X"00000000",
		16#0364# => X"00000000",
		16#0365# => X"00000000",
		16#0366# => X"00000000",
		16#0367# => X"00000000",
		16#0368# => X"00000000",
		16#0369# => X"00000000",
		16#036a# => X"00000000",
		16#036b# => X"00000000",
		16#036c# => X"00000000",
		16#036d# => X"00000000",
		16#036e# => X"00000000",
		16#036f# => X"00000000",
		16#0370# => X"00000000",
		16#0371# => X"00000000",
		16#0372# => X"00000000",
		16#0373# => X"00000000",
		16#0374# => X"00000000",
		16#0375# => X"00000000",
		16#0376# => X"00000000",
		16#0377# => X"00000000",
		16#0378# => X"00000000",
		16#0379# => X"00000000",
		16#037a# => X"00000000",
		16#037b# => X"00000000",
		16#037c# => X"00000000",
		16#037d# => X"00000000",
		16#037e# => X"00000000",
		16#037f# => X"00000000",
		16#0380# => X"00000000",
		16#0381# => X"00000000",
		16#0382# => X"00000000",
		16#0383# => X"00000000",
		16#0384# => X"00000000",
		16#0385# => X"00000000",
		16#0386# => X"00000000",
		16#0387# => X"00000000",
		16#0388# => X"00000000",
		16#0389# => X"00000000",
		16#038a# => X"00000000",
		16#038b# => X"00000000",
		16#038c# => X"00000000",
		16#038d# => X"00000000",
		16#038e# => X"00000000",
		16#038f# => X"00000000",
		16#0390# => X"00000000",
		16#0391# => X"00000000",
		16#0392# => X"00000000",
		16#0393# => X"00000000",
		16#0394# => X"00000000",
		16#0395# => X"00000000",
		16#0396# => X"00000000",
		16#0397# => X"00000000",
		16#0398# => X"00000000",
		16#0399# => X"00000000",
		16#039a# => X"00000000",
		16#039b# => X"00000000",
		16#039c# => X"00000000",
		16#039d# => X"00000000",
		16#039e# => X"00000000",
		16#039f# => X"00000000",
		16#03a0# => X"00000000",
		16#03a1# => X"00000000",
		16#03a2# => X"00000000",
		16#03a3# => X"00000000",
		16#03a4# => X"00000000",
		16#03a5# => X"00000000",
		16#03a6# => X"00000000",
		16#03a7# => X"00000000",
		16#03a8# => X"00000000",
		16#03a9# => X"00000000",
		16#03aa# => X"00000000",
		16#03ab# => X"00000000",
		16#03ac# => X"00000000",
		16#03ad# => X"00000000",
		16#03ae# => X"00000000",
		16#03af# => X"00000000",
		16#03b0# => X"00000000",
		16#03b1# => X"00000000",
		16#03b2# => X"00000000",
		16#03b3# => X"00000000",
		16#03b4# => X"00000000",
		16#03b5# => X"00000000",
		16#03b6# => X"00000000",
		16#03b7# => X"00000000",
		16#03b8# => X"00000000",
		16#03b9# => X"00000000",
		16#03ba# => X"00000000",
		16#03bb# => X"00000000",
		16#03bc# => X"00000000",
		16#03bd# => X"00000000",
		16#03be# => X"00000000",
		16#03bf# => X"00000000",
		16#03c0# => X"00000000",
		16#03c1# => X"00000000",
		16#03c2# => X"00000000",
		16#03c3# => X"00000000",
		16#03c4# => X"00000000",
		16#03c5# => X"00000000",
		16#03c6# => X"00000000",
		16#03c7# => X"00000000",
		16#03c8# => X"00000000",
		16#03c9# => X"00000000",
		16#03ca# => X"00000000",
		16#03cb# => X"00000000",
		16#03cc# => X"00000000",
		16#03cd# => X"00000000",
		16#03ce# => X"00000000",
		16#03cf# => X"00000000",
		16#03d0# => X"00000000",
		16#03d1# => X"00000000",
		16#03d2# => X"00000000",
		16#03d3# => X"00000000",
		16#03d4# => X"00000000",
		16#03d5# => X"00000000",
		16#03d6# => X"00000000",
		16#03d7# => X"00000000",
		16#03d8# => X"00000000",
		16#03d9# => X"00000000",
		16#03da# => X"00000000",
		16#03db# => X"00000000",
		16#03dc# => X"00000000",
		16#03dd# => X"00000000",
		16#03de# => X"00000000",
		16#03df# => X"00000000",
		16#03e0# => X"00000000",
		16#03e1# => X"00000000",
		16#03e2# => X"00000000",
		16#03e3# => X"00000000",
		16#03e4# => X"00000000",
		16#03e5# => X"00000000",
		16#03e6# => X"00000000",
		16#03e7# => X"00000000",
		16#03e8# => X"00000000",
		16#03e9# => X"00000000",
		16#03ea# => X"00000000",
		16#03eb# => X"00000000",
		16#03ec# => X"00000000",
		16#03ed# => X"00000000",
		16#03ee# => X"00000000",
		16#03ef# => X"00000000",
		16#03f0# => X"00000000",
		16#03f1# => X"00000000",
		16#03f2# => X"00000000",
		16#03f3# => X"00000000",
		16#03f4# => X"00000000",
		16#03f5# => X"00000000",
		16#03f6# => X"00000000",
		16#03f7# => X"00000000",
		16#03f8# => X"00000000",
		16#03f9# => X"00000000",
		16#03fa# => X"00000000",
		16#03fb# => X"00000000",
		16#03fc# => X"00000000",
		16#03fd# => X"00000000",
		16#03fe# => X"00000000",
		16#03ff# => X"00000000",
		16#0400# => X"00000000",
		16#0401# => X"00000000",
		16#0402# => X"00000000",
		16#0403# => X"00000000",
		16#0404# => X"00000000",
		16#0405# => X"00000000",
		16#0406# => X"00000000",
		16#0407# => X"00000000",
		16#0408# => X"00000000",
		16#0409# => X"00000000",
		16#040a# => X"00000000",
		16#040b# => X"00000000",
		16#040c# => X"00000000",
		16#040d# => X"00000000",
		16#040e# => X"00000000",
		16#040f# => X"00000000",
		16#0410# => X"00000000",
		16#0411# => X"00000000",
		16#0412# => X"13052500",
		16#0413# => X"b305b500",
		16#0414# => X"2320b600",
		16#0415# => X"67800000",
		16#0416# => X"130101fe",
		16#0417# => X"23263101",
		16#0418# => X"93095600",
		16#0419# => X"232a9100",
		16#041a# => X"93942900",
		16#041b# => X"232c8100",
		16#041c# => X"23282101",
		16#041d# => X"232e1100",
		16#041e# => X"b3049500",
		16#041f# => X"13090600",
		16#0420# => X"13840500",
		16#0421# => X"23ac3407",
		16#0422# => X"23a0d400",
		16#0423# => X"23a2d400",
		16#0424# => X"13850900",
		16#0425# => X"9305800c",
		16#0426# => X"ef108159",
		16#0427# => X"13192900",
		16#0428# => X"b3072501",
		16#0429# => X"b307f400",
		16#042a# => X"03a70701",
		16#042b# => X"23aa3701",
		16#042c# => X"23ac3701",
		16#042d# => X"13071700",
		16#042e# => X"23a8e700",
		16#042f# => X"83a70400",
		16#0430# => X"3304a400",
		16#0431# => X"33042401",
		16#0432# => X"37160000",
		16#0433# => X"33048600",
		16#0434# => X"232af4fa",
		16#0435# => X"8320c101",
		16#0436# => X"03248101",
		16#0437# => X"b7870110",
		16#0438# => X"13075000",
		16#0439# => X"23a4e79c",
		16#043a# => X"83244101",
		16#043b# => X"03290101",
		16#043c# => X"8329c100",
		16#043d# => X"13010102",
		16#043e# => X"67800000",
		16#043f# => X"1375f50f",
		16#0440# => X"93f5f50f",
		16#0441# => X"6306b500",
		16#0442# => X"13050000",
		16#0443# => X"67800000",
		16#0444# => X"b7870110",
		16#0445# => X"2386a79c",
		16#0446# => X"13051000",
		16#0447# => X"67800000",
		16#0448# => X"130101ff",
		16#0449# => X"23248100",
		16#044a# => X"23229100",
		16#044b# => X"23261100",
		16#044c# => X"13040500",
		16#044d# => X"93840500",
		16#044e# => X"83c53400",
		16#044f# => X"03452400",
		16#0450# => X"eff0dffb",
		16#0451# => X"e31a05fe",
		16#0452# => X"93850400",
		16#0453# => X"13050400",
		16#0454# => X"ef008054",
		16#0455# => X"93070000",
		16#0456# => X"635aa000",
		16#0457# => X"b7870110",
		16#0458# => X"1307a000",
		16#0459# => X"23a4e79c",
		16#045a# => X"93071000",
		16#045b# => X"8320c100",
		16#045c# => X"03248100",
		16#045d# => X"83244100",
		16#045e# => X"13850700",
		16#045f# => X"13010101",
		16#0460# => X"67800000",
		16#0461# => X"1305e5ff",
		16#0462# => X"13351500",
		16#0463# => X"67800000",
		16#0464# => X"130101ff",
		16#0465# => X"23248100",
		16#0466# => X"23229100",
		16#0467# => X"23261100",
		16#0468# => X"13040500",
		16#0469# => X"93840500",
		16#046a# => X"eff0dffd",
		16#046b# => X"630e0502",
		16#046c# => X"23a08400",
		16#046d# => X"93071000",
		16#046e# => X"6300f404",
		16#046f# => X"63060404",
		16#0470# => X"13072000",
		16#0471# => X"630ee404",
		16#0472# => X"93074000",
		16#0473# => X"6314f400",
		16#0474# => X"23a0e400",
		16#0475# => X"8320c100",
		16#0476# => X"03248100",
		16#0477# => X"83244100",
		16#0478# => X"13010101",
		16#0479# => X"67800000",
		16#047a# => X"93073000",
		16#047b# => X"23a0f400",
		16#047c# => X"93071000",
		16#047d# => X"e314f4fc",
		16#047e# => X"b7870110",
		16#047f# => X"03a7879c",
		16#0480# => X"93074006",
		16#0481# => X"63dae702",
		16#0482# => X"8320c100",
		16#0483# => X"03248100",
		16#0484# => X"23a00400",
		16#0485# => X"83244100",
		16#0486# => X"13010101",
		16#0487# => X"67800000",
		16#0488# => X"8320c100",
		16#0489# => X"03248100",
		16#048a# => X"23a0f400",
		16#048b# => X"83244100",
		16#048c# => X"13010101",
		16#048d# => X"67800000",
		16#048e# => X"8320c100",
		16#048f# => X"03248100",
		16#0490# => X"93073000",
		16#0491# => X"23a0f400",
		16#0492# => X"83244100",
		16#0493# => X"13010101",
		16#0494# => X"67800000",
		16#0495# => X"130101fe",
		16#0496# => X"2322b100",
		16#0497# => X"2324c100",
		16#0498# => X"2326d100",
		16#0499# => X"2328e100",
		16#049a# => X"232af100",
		16#049b# => X"232c0101",
		16#049c# => X"232e1101",
		16#049d# => X"13010102",
		16#049e# => X"67800000",
		16#049f# => X"b7870110",
		16#04a0# => X"03c7c79c",
		16#04a1# => X"93071004",
		16#04a2# => X"6304f700",
		16#04a3# => X"67800000",
		16#04a4# => X"83270500",
		16#04a5# => X"37870110",
		16#04a6# => X"0327879c",
		16#04a7# => X"93879700",
		16#04a8# => X"b387e740",
		16#04a9# => X"2320f500",
		16#04aa# => X"67800000",
		16#04ab# => X"b7870110",
		16#04ac# => X"03a6079d",
		16#04ad# => X"63080600",
		16#04ae# => X"03270600",
		16#04af# => X"2320e500",
		16#04b0# => X"03a6079d",
		16#04b1# => X"b7870110",
		16#04b2# => X"83a5879c",
		16#04b3# => X"1306c600",
		16#04b4# => X"1305a000",
		16#04b5# => X"6ff05fd7",
		16#04b6# => X"130101ff",
		16#04b7# => X"23202101",
		16#04b8# => X"37890110",
		16#04b9# => X"8327099d",
		16#04ba# => X"23248100",
		16#04bb# => X"03240500",
		16#04bc# => X"03a70700",
		16#04bd# => X"23229100",
		16#04be# => X"83ae4700",
		16#04bf# => X"03ae8700",
		16#04c0# => X"03a30701",
		16#04c1# => X"83a84701",
		16#04c2# => X"03a88701",
		16#04c3# => X"83a50702",
		16#04c4# => X"03a64702",
		16#04c5# => X"83a68702",
		16#04c6# => X"23261100",
		16#04c7# => X"93040500",
		16#04c8# => X"03a5c701",
		16#04c9# => X"83a7c702",
		16#04ca# => X"2320e400",
		16#04cb# => X"03a70400",
		16#04cc# => X"232ea400",
		16#04cd# => X"2326f402",
		16#04ce# => X"2322d401",
		16#04cf# => X"93075000",
		16#04d0# => X"2324c401",
		16#04d1# => X"23286400",
		16#04d2# => X"232a1401",
		16#04d3# => X"232c0401",
		16#04d4# => X"2320b402",
		16#04d5# => X"2322c402",
		16#04d6# => X"2324d402",
		16#04d7# => X"23a6f400",
		16#04d8# => X"2326f400",
		16#04d9# => X"2320e400",
		16#04da# => X"13050400",
		16#04db# => X"eff01ff4",
		16#04dc# => X"83274400",
		16#04dd# => X"63800708",
		16#04de# => X"83a70400",
		16#04df# => X"8320c100",
		16#04e0# => X"03248100",
		16#04e1# => X"83af0700",
		16#04e2# => X"03af4700",
		16#04e3# => X"83ae8700",
		16#04e4# => X"03aec700",
		16#04e5# => X"03a30701",
		16#04e6# => X"83a84701",
		16#04e7# => X"03a88701",
		16#04e8# => X"83a5c701",
		16#04e9# => X"03a60702",
		16#04ea# => X"83a64702",
		16#04eb# => X"03a78702",
		16#04ec# => X"83a7c702",
		16#04ed# => X"23a0f401",
		16#04ee# => X"23a2e401",
		16#04ef# => X"23a4d401",
		16#04f0# => X"23a6c401",
		16#04f1# => X"23a86400",
		16#04f2# => X"23aa1401",
		16#04f3# => X"23ac0401",
		16#04f4# => X"23aeb400",
		16#04f5# => X"23a0c402",
		16#04f6# => X"23a2d402",
		16#04f7# => X"23a4e402",
		16#04f8# => X"23a6f402",
		16#04f9# => X"03290100",
		16#04fa# => X"83244100",
		16#04fb# => X"13010101",
		16#04fc# => X"67800000",
		16#04fd# => X"03a58400",
		16#04fe# => X"93076000",
		16#04ff# => X"93058400",
		16#0500# => X"2326f400",
		16#0501# => X"eff0dfd8",
		16#0502# => X"8327099d",
		16#0503# => X"0325c400",
		16#0504# => X"1306c400",
		16#0505# => X"83a70700",
		16#0506# => X"8320c100",
		16#0507# => X"83244100",
		16#0508# => X"2320f400",
		16#0509# => X"03248100",
		16#050a# => X"03290100",
		16#050b# => X"9305a000",
		16#050c# => X"13010101",
		16#050d# => X"6ff05fc1",
		16#050e# => X"b7870110",
		16#050f# => X"83c7c79c",
		16#0510# => X"37870110",
		16#0511# => X"832607aa",
		16#0512# => X"9387f7fb",
		16#0513# => X"93b71700",
		16#0514# => X"b3e7d700",
		16#0515# => X"2320f7aa",
		16#0516# => X"b7870110",
		16#0517# => X"13072004",
		16#0518# => X"a386e79c",
		16#0519# => X"67800000",
		16#051a# => X"b7870110",
		16#051b# => X"13071004",
		16#051c# => X"2386e79c",
		16#051d# => X"b7870110",
		16#051e# => X"23a007aa",
		16#051f# => X"67800000",
		16#0520# => X"130101fc",
		16#0521# => X"2324c102",
		16#0522# => X"2326d102",
		16#0523# => X"2328e102",
		16#0524# => X"232af102",
		16#0525# => X"232c0103",
		16#0526# => X"232e1103",
		16#0527# => X"13860500",
		16#0528# => X"83258500",
		16#0529# => X"93068102",
		16#052a# => X"232e1100",
		16#052b# => X"2326d100",
		16#052c# => X"ef004039",
		16#052d# => X"8320c101",
		16#052e# => X"13010104",
		16#052f# => X"67800000",
		16#0530# => X"130101fc",
		16#0531# => X"232af102",
		16#0532# => X"83a7c181",
		16#0533# => X"2324c102",
		16#0534# => X"2326d102",
		16#0535# => X"2322b102",
		16#0536# => X"2328e102",
		16#0537# => X"232c0103",
		16#0538# => X"232e1103",
		16#0539# => X"83a58700",
		16#053a# => X"93064102",
		16#053b# => X"13060500",
		16#053c# => X"13850700",
		16#053d# => X"232e1100",
		16#053e# => X"2326d100",
		16#053f# => X"ef008034",
		16#0540# => X"8320c101",
		16#0541# => X"13010104",
		16#0542# => X"67800000",
		16#0543# => X"03268500",
		16#0544# => X"6f008001",
		16#0545# => X"83a7c181",
		16#0546# => X"93050500",
		16#0547# => X"03a68700",
		16#0548# => X"13850700",
		16#0549# => X"6f004000",
		16#054a# => X"130101fe",
		16#054b# => X"232c8100",
		16#054c# => X"232e1100",
		16#054d# => X"13040500",
		16#054e# => X"63000502",
		16#054f# => X"83278503",
		16#0550# => X"639c0700",
		16#0551# => X"2326c100",
		16#0552# => X"2324b100",
		16#0553# => X"ef20d019",
		16#0554# => X"0326c100",
		16#0555# => X"83258100",
		16#0556# => X"83278600",
		16#0557# => X"9387f7ff",
		16#0558# => X"2324f600",
		16#0559# => X"63d60702",
		16#055a# => X"03278601",
		16#055b# => X"63c8e700",
		16#055c# => X"93f7f50f",
		16#055d# => X"1307a000",
		16#055e# => X"639ce700",
		16#055f# => X"13050400",
		16#0560# => X"03248101",
		16#0561# => X"8320c101",
		16#0562# => X"13010102",
		16#0563# => X"6f204034",
		16#0564# => X"83270600",
		16#0565# => X"13f5f50f",
		16#0566# => X"13871700",
		16#0567# => X"2320e600",
		16#0568# => X"2380b700",
		16#0569# => X"8320c101",
		16#056a# => X"03248101",
		16#056b# => X"13010102",
		16#056c# => X"67800000",
		16#056d# => X"13860500",
		16#056e# => X"93050500",
		16#056f# => X"03a5c181",
		16#0570# => X"6ff09ff6",
		16#0571# => X"130101fc",
		16#0572# => X"232c8102",
		16#0573# => X"13040500",
		16#0574# => X"13850500",
		16#0575# => X"2326b100",
		16#0576# => X"232e1102",
		16#0577# => X"ef008023",
		16#0578# => X"b7470110",
		16#0579# => X"9387c79d",
		16#057a# => X"2324f102",
		16#057b# => X"93071000",
		16#057c# => X"2326f102",
		16#057d# => X"93070102",
		16#057e# => X"8325c100",
		16#057f# => X"232af100",
		16#0580# => X"93072000",
		16#0581# => X"232cf100",
		16#0582# => X"83278403",
		16#0583# => X"2322a102",
		16#0584# => X"13051500",
		16#0585# => X"2320b102",
		16#0586# => X"232ea100",
		16#0587# => X"83258400",
		16#0588# => X"639a0700",
		16#0589# => X"13050400",
		16#058a# => X"2326b100",
		16#058b# => X"ef20d00b",
		16#058c# => X"8325c100",
		16#058d# => X"8397c500",
		16#058e# => X"13972701",
		16#058f# => X"63420702",
		16#0590# => X"b7260000",
		16#0591# => X"03a74506",
		16#0592# => X"b3e7d700",
		16#0593# => X"2396f500",
		16#0594# => X"b7e7ffff",
		16#0595# => X"9387f7ff",
		16#0596# => X"b377f700",
		16#0597# => X"23a2f506",
		16#0598# => X"13064101",
		16#0599# => X"13050400",
		16#059a# => X"ef201059",
		16#059b# => X"9307f0ff",
		16#059c# => X"63140500",
		16#059d# => X"9307a000",
		16#059e# => X"8320c103",
		16#059f# => X"03248103",
		16#05a0# => X"13850700",
		16#05a1# => X"13010104",
		16#05a2# => X"67800000",
		16#05a3# => X"93050500",
		16#05a4# => X"03a5c181",
		16#05a5# => X"6ff01ff3",
		16#05a6# => X"3367b500",
		16#05a7# => X"9303f0ff",
		16#05a8# => X"13773700",
		16#05a9# => X"63100710",
		16#05aa# => X"b7877f7f",
		16#05ab# => X"9387f7f7",
		16#05ac# => X"03260500",
		16#05ad# => X"83a60500",
		16#05ae# => X"b372f600",
		16#05af# => X"3363f600",
		16#05b0# => X"b382f200",
		16#05b1# => X"b3e26200",
		16#05b2# => X"63927210",
		16#05b3# => X"6316d608",
		16#05b4# => X"03264500",
		16#05b5# => X"83a64500",
		16#05b6# => X"b372f600",
		16#05b7# => X"3363f600",
		16#05b8# => X"b382f200",
		16#05b9# => X"b3e26200",
		16#05ba# => X"639e720c",
		16#05bb# => X"6316d606",
		16#05bc# => X"03268500",
		16#05bd# => X"83a68500",
		16#05be# => X"b372f600",
		16#05bf# => X"3363f600",
		16#05c0# => X"b382f200",
		16#05c1# => X"b3e26200",
		16#05c2# => X"6398720c",
		16#05c3# => X"6316d604",
		16#05c4# => X"0326c500",
		16#05c5# => X"83a6c500",
		16#05c6# => X"b372f600",
		16#05c7# => X"3363f600",
		16#05c8# => X"b382f200",
		16#05c9# => X"b3e26200",
		16#05ca# => X"6392720c",
		16#05cb# => X"6316d602",
		16#05cc# => X"03260501",
		16#05cd# => X"83a60501",
		16#05ce# => X"b372f600",
		16#05cf# => X"3363f600",
		16#05d0# => X"b382f200",
		16#05d1# => X"b3e26200",
		16#05d2# => X"639c720a",
		16#05d3# => X"13054501",
		16#05d4# => X"93854501",
		16#05d5# => X"e30ed6f4",
		16#05d6# => X"13170601",
		16#05d7# => X"93970601",
		16#05d8# => X"631ef700",
		16#05d9# => X"13570601",
		16#05da# => X"93d70601",
		16#05db# => X"3305f740",
		16#05dc# => X"9375f50f",
		16#05dd# => X"63900502",
		16#05de# => X"67800000",
		16#05df# => X"13570701",
		16#05e0# => X"93d70701",
		16#05e1# => X"3305f740",
		16#05e2# => X"9375f50f",
		16#05e3# => X"63940500",
		16#05e4# => X"67800000",
		16#05e5# => X"1377f70f",
		16#05e6# => X"93f7f70f",
		16#05e7# => X"3305f740",
		16#05e8# => X"67800000",
		16#05e9# => X"03460500",
		16#05ea# => X"83c60500",
		16#05eb# => X"13051500",
		16#05ec# => X"93851500",
		16#05ed# => X"6314d600",
		16#05ee# => X"e31606fe",
		16#05ef# => X"3305d640",
		16#05f0# => X"67800000",
		16#05f1# => X"13054500",
		16#05f2# => X"93854500",
		16#05f3# => X"e31cd6fc",
		16#05f4# => X"13050000",
		16#05f5# => X"67800000",
		16#05f6# => X"13058500",
		16#05f7# => X"93858500",
		16#05f8# => X"e312d6fc",
		16#05f9# => X"13050000",
		16#05fa# => X"67800000",
		16#05fb# => X"1305c500",
		16#05fc# => X"9385c500",
		16#05fd# => X"e318d6fa",
		16#05fe# => X"13050000",
		16#05ff# => X"67800000",
		16#0600# => X"13050501",
		16#0601# => X"93850501",
		16#0602# => X"e31ed6f8",
		16#0603# => X"13050000",
		16#0604# => X"67800000",
		16#0605# => X"93070500",
		16#0606# => X"93871700",
		16#0607# => X"03c7f7ff",
		16#0608# => X"e31c07fe",
		16#0609# => X"3385a740",
		16#060a# => X"1305f5ff",
		16#060b# => X"67800000",
		16#060c# => X"93050500",
		16#060d# => X"03a5c181",
		16#060e# => X"6f004000",
		16#060f# => X"13850500",
		16#0610# => X"6fb0905c",
		16#0611# => X"130101e2",
		16#0612# => X"232e111c",
		16#0613# => X"232a911c",
		16#0614# => X"2328211d",
		16#0615# => X"2326311d",
		16#0616# => X"232c811b",
		16#0617# => X"13890500",
		16#0618# => X"93040600",
		16#0619# => X"138c0600",
		16#061a# => X"232c811c",
		16#061b# => X"2324411d",
		16#061c# => X"2322511d",
		16#061d# => X"2320611d",
		16#061e# => X"232e711b",
		16#061f# => X"232a911b",
		16#0620# => X"2328a11b",
		16#0621# => X"2326b11b",
		16#0622# => X"93090500",
		16#0623# => X"ef50401a",
		16#0624# => X"83270500",
		16#0625# => X"13850700",
		16#0626# => X"232cf102",
		16#0627# => X"eff09ff7",
		16#0628# => X"2322a102",
		16#0629# => X"2320010e",
		16#062a# => X"2322010e",
		16#062b# => X"2324010e",
		16#062c# => X"2326010e",
		16#062d# => X"638a0900",
		16#062e# => X"83a78903",
		16#062f# => X"63960700",
		16#0630# => X"13850900",
		16#0631# => X"ef204062",
		16#0632# => X"8317c900",
		16#0633# => X"13972701",
		16#0634# => X"63420702",
		16#0635# => X"b7260000",
		16#0636# => X"03274906",
		16#0637# => X"b3e7d700",
		16#0638# => X"2316f900",
		16#0639# => X"b7e7ffff",
		16#063a# => X"9387f7ff",
		16#063b# => X"b377f700",
		16#063c# => X"2322f906",
		16#063d# => X"8357c900",
		16#063e# => X"93f78700",
		16#063f# => X"638e0706",
		16#0640# => X"83270901",
		16#0641# => X"638a0706",
		16#0642# => X"8357c900",
		16#0643# => X"1307a000",
		16#0644# => X"93f7a701",
		16#0645# => X"6390e708",
		16#0646# => X"8317e900",
		16#0647# => X"63cc0706",
		16#0648# => X"93060c00",
		16#0649# => X"13860400",
		16#064a# => X"93050900",
		16#064b# => X"13850900",
		16#064c# => X"ef10506e",
		16#064d# => X"2324a102",
		16#064e# => X"8320c11d",
		16#064f# => X"0324811d",
		16#0650# => X"03258102",
		16#0651# => X"8324411d",
		16#0652# => X"0329011d",
		16#0653# => X"8329c11c",
		16#0654# => X"032a811c",
		16#0655# => X"832a411c",
		16#0656# => X"032b011c",
		16#0657# => X"832bc11b",
		16#0658# => X"032c811b",
		16#0659# => X"832c411b",
		16#065a# => X"032d011b",
		16#065b# => X"832dc11a",
		16#065c# => X"1301011e",
		16#065d# => X"67800000",
		16#065e# => X"93050900",
		16#065f# => X"13850900",
		16#0660# => X"ef200009",
		16#0661# => X"e30205f8",
		16#0662# => X"9307f0ff",
		16#0663# => X"2324f102",
		16#0664# => X"6ff09ffa",
		16#0665# => X"b7470110",
		16#0666# => X"938787b5",
		16#0667# => X"2328f104",
		16#0668# => X"b7470110",
		16#0669# => X"9308c10f",
		16#066a# => X"938747cd",
		16#066b# => X"232a110d",
		16#066c# => X"232e010c",
		16#066d# => X"232c010c",
		16#066e# => X"130a0000",
		16#066f# => X"138d0800",
		16#0670# => X"23220104",
		16#0671# => X"23200104",
		16#0672# => X"232a0100",
		16#0673# => X"232a0102",
		16#0674# => X"232e0102",
		16#0675# => X"23240102",
		16#0676# => X"232cf100",
		16#0677# => X"13840400",
		16#0678# => X"13075002",
		16#0679# => X"83470400",
		16#067a# => X"63840700",
		16#067b# => X"6392e70c",
		16#067c# => X"b30a9440",
		16#067d# => X"638a0a04",
		16#067e# => X"8327c10d",
		16#067f# => X"23209d00",
		16#0680# => X"23225d01",
		16#0681# => X"b3875701",
		16#0682# => X"232ef10c",
		16#0683# => X"8327810d",
		16#0684# => X"13077000",
		16#0685# => X"130d8d00",
		16#0686# => X"93871700",
		16#0687# => X"232cf10c",
		16#0688# => X"635ef700",
		16#0689# => X"1306410d",
		16#068a# => X"93050900",
		16#068b# => X"13850900",
		16#068c# => X"ef908032",
		16#068d# => X"63180578",
		16#068e# => X"130dc10f",
		16#068f# => X"83278102",
		16#0690# => X"b3875701",
		16#0691# => X"2324f102",
		16#0692# => X"83470400",
		16#0693# => X"63940700",
		16#0694# => X"6f101059",
		16#0695# => X"93071400",
		16#0696# => X"2320f102",
		16#0697# => X"a30b010a",
		16#0698# => X"130bf0ff",
		16#0699# => X"23260102",
		16#069a# => X"13040000",
		16#069b# => X"930a9000",
		16#069c# => X"930ba005",
		16#069d# => X"83270102",
		16#069e# => X"83c70700",
		16#069f# => X"2326f100",
		16#06a0# => X"83270102",
		16#06a1# => X"93871700",
		16#06a2# => X"2320f102",
		16#06a3# => X"8327c100",
		16#06a4# => X"938707fe",
		16#06a5# => X"63f4fb00",
		16#06a6# => X"6f10c024",
		16#06a7# => X"03270105",
		16#06a8# => X"93972700",
		16#06a9# => X"b387e700",
		16#06aa# => X"83a70700",
		16#06ab# => X"67800700",
		16#06ac# => X"13041400",
		16#06ad# => X"6ff01ff3",
		16#06ae# => X"b7470110",
		16#06af# => X"93878791",
		16#06b0# => X"2322f104",
		16#06b1# => X"93770402",
		16#06b2# => X"63940700",
		16#06b3# => X"6f10c004",
		16#06b4# => X"130c7c00",
		16#06b5# => X"137c8cff",
		16#06b6# => X"93078c00",
		16#06b7# => X"832c0c00",
		16#06b8# => X"032c4c00",
		16#06b9# => X"232ef100",
		16#06ba# => X"93771400",
		16#06bb# => X"63800702",
		16#06bc# => X"b3e78c01",
		16#06bd# => X"638c0700",
		16#06be# => X"93070003",
		16#06bf# => X"230cf10a",
		16#06c0# => X"8347c100",
		16#06c1# => X"13642400",
		16#06c2# => X"a30cf10a",
		16#06c3# => X"1374f4bf",
		16#06c4# => X"93072000",
		16#06c5# => X"6f00106a",
		16#06c6# => X"13850900",
		16#06c7# => X"ef405071",
		16#06c8# => X"83274500",
		16#06c9# => X"13850700",
		16#06ca# => X"232ef102",
		16#06cb# => X"eff09fce",
		16#06cc# => X"232aa102",
		16#06cd# => X"13850900",
		16#06ce# => X"ef40906f",
		16#06cf# => X"83278500",
		16#06d0# => X"232af100",
		16#06d1# => X"83274103",
		16#06d2# => X"e38407f2",
		16#06d3# => X"83274101",
		16#06d4# => X"e38007f2",
		16#06d5# => X"83c70700",
		16#06d6# => X"e38c07f0",
		16#06d7# => X"13640440",
		16#06d8# => X"6ff01ff1",
		16#06d9# => X"8347710b",
		16#06da# => X"e39407f0",
		16#06db# => X"93070002",
		16#06dc# => X"a30bf10a",
		16#06dd# => X"6ff0dfef",
		16#06de# => X"13641400",
		16#06df# => X"6ff05fef",
		16#06e0# => X"83270c00",
		16#06e1# => X"130c4c00",
		16#06e2# => X"2326f102",
		16#06e3# => X"e3d207ee",
		16#06e4# => X"b307f040",
		16#06e5# => X"2326f102",
		16#06e6# => X"13644400",
		16#06e7# => X"6ff05fed",
		16#06e8# => X"9307b002",
		16#06e9# => X"6ff0dffc",
		16#06ea# => X"83270102",
		16#06eb# => X"1307a002",
		16#06ec# => X"938c1700",
		16#06ed# => X"83c70700",
		16#06ee# => X"2326f100",
		16#06ef# => X"6398e704",
		16#06f0# => X"032b0c00",
		16#06f1# => X"93074c00",
		16#06f2# => X"63540b00",
		16#06f3# => X"130bf0ff",
		16#06f4# => X"138c0700",
		16#06f5# => X"23209103",
		16#06f6# => X"6ff09fe9",
		16#06f7# => X"13050b00",
		16#06f8# => X"9305a000",
		16#06f9# => X"ef00d124",
		16#06fa# => X"938c1c00",
		16#06fb# => X"83c7fcff",
		16#06fc# => X"330bb501",
		16#06fd# => X"2326f100",
		16#06fe# => X"8327c100",
		16#06ff# => X"938d07fd",
		16#0700# => X"e3febafd",
		16#0701# => X"23209103",
		16#0702# => X"6ff05fe8",
		16#0703# => X"130b0000",
		16#0704# => X"6ff09ffe",
		16#0705# => X"13640408",
		16#0706# => X"6ff09fe5",
		16#0707# => X"832c0102",
		16#0708# => X"23260102",
		16#0709# => X"0325c102",
		16#070a# => X"9305a000",
		16#070b# => X"938c1c00",
		16#070c# => X"ef001120",
		16#070d# => X"8327c100",
		16#070e# => X"938707fd",
		16#070f# => X"b387a700",
		16#0710# => X"2326f102",
		16#0711# => X"83c7fcff",
		16#0712# => X"2326f100",
		16#0713# => X"938707fd",
		16#0714# => X"e3fafafc",
		16#0715# => X"6ff01ffb",
		16#0716# => X"13648400",
		16#0717# => X"6ff05fe1",
		16#0718# => X"83270102",
		16#0719# => X"03c70700",
		16#071a# => X"93078006",
		16#071b# => X"631cf700",
		16#071c# => X"83270102",
		16#071d# => X"13640420",
		16#071e# => X"93871700",
		16#071f# => X"2320f102",
		16#0720# => X"6ff01fdf",
		16#0721# => X"13640404",
		16#0722# => X"6ff09fde",
		16#0723# => X"83270102",
		16#0724# => X"03c70700",
		16#0725# => X"9307c006",
		16#0726# => X"631cf700",
		16#0727# => X"83270102",
		16#0728# => X"93871700",
		16#0729# => X"2320f102",
		16#072a# => X"13640402",
		16#072b# => X"6ff05fdc",
		16#072c# => X"13640401",
		16#072d# => X"6ff0dfdb",
		16#072e# => X"93074c00",
		16#072f# => X"232ef100",
		16#0730# => X"83270c00",
		16#0731# => X"a30b010a",
		16#0732# => X"230ef112",
		16#0733# => X"23280100",
		16#0734# => X"130b1000",
		16#0735# => X"930a0000",
		16#0736# => X"130c0000",
		16#0737# => X"930b0000",
		16#0738# => X"930c0000",
		16#0739# => X"9304c113",
		16#073a# => X"23285103",
		16#073b# => X"63d46a01",
		16#073c# => X"23286103",
		16#073d# => X"0347710b",
		16#073e# => X"63080700",
		16#073f# => X"83270103",
		16#0740# => X"93871700",
		16#0741# => X"2328f102",
		16#0742# => X"937d2400",
		16#0743# => X"63880d00",
		16#0744# => X"83270103",
		16#0745# => X"93872700",
		16#0746# => X"2328f102",
		16#0747# => X"93774408",
		16#0748# => X"2324f104",
		16#0749# => X"639c0706",
		16#074a# => X"8327c102",
		16#074b# => X"03270103",
		16#074c# => X"3387e740",
		16#074d# => X"6354e006",
		16#074e# => X"374e0110",
		16#074f# => X"930e0001",
		16#0750# => X"130e4ecc",
		16#0751# => X"130f7000",
		16#0752# => X"8326810d",
		16#0753# => X"2320cd01",
		16#0754# => X"0326c10d",
		16#0755# => X"93861600",
		16#0756# => X"93058d00",
		16#0757# => X"63d4ee00",
		16#0758# => X"6f00107a",
		16#0759# => X"2322ed00",
		16#075a# => X"3307c700",
		16#075b# => X"232ee10c",
		16#075c# => X"232cd10c",
		16#075d# => X"13077000",
		16#075e# => X"138d0500",
		16#075f# => X"6350d702",
		16#0760# => X"1306410d",
		16#0761# => X"93050900",
		16#0762# => X"13850900",
		16#0763# => X"ef80d07c",
		16#0764# => X"63040500",
		16#0765# => X"6f10901e",
		16#0766# => X"130dc10f",
		16#0767# => X"0347710b",
		16#0768# => X"630a0704",
		16#0769# => X"1307710b",
		16#076a# => X"2320ed00",
		16#076b# => X"13071000",
		16#076c# => X"2322ed00",
		16#076d# => X"0327c10d",
		16#076e# => X"93067000",
		16#076f# => X"130d8d00",
		16#0770# => X"13071700",
		16#0771# => X"232ee10c",
		16#0772# => X"0327810d",
		16#0773# => X"13071700",
		16#0774# => X"232ce10c",
		16#0775# => X"63d0e602",
		16#0776# => X"1306410d",
		16#0777# => X"93050900",
		16#0778# => X"13850900",
		16#0779# => X"ef805077",
		16#077a# => X"63040500",
		16#077b# => X"6f101019",
		16#077c# => X"130dc10f",
		16#077d# => X"638a0d04",
		16#077e# => X"1307810b",
		16#077f# => X"2320ed00",
		16#0780# => X"13072000",
		16#0781# => X"2322ed00",
		16#0782# => X"0327c10d",
		16#0783# => X"93067000",
		16#0784# => X"130d8d00",
		16#0785# => X"13072700",
		16#0786# => X"232ee10c",
		16#0787# => X"0327810d",
		16#0788# => X"13071700",
		16#0789# => X"232ce10c",
		16#078a# => X"63d0e602",
		16#078b# => X"1306410d",
		16#078c# => X"93050900",
		16#078d# => X"13850900",
		16#078e# => X"ef801072",
		16#078f# => X"63040500",
		16#0790# => X"6f10d013",
		16#0791# => X"130dc10f",
		16#0792# => X"83278104",
		16#0793# => X"13070008",
		16#0794# => X"6398e706",
		16#0795# => X"8327c102",
		16#0796# => X"03270103",
		16#0797# => X"b38de740",
		16#0798# => X"6350b007",
		16#0799# => X"93070001",
		16#079a# => X"130e7000",
		16#079b# => X"0327810d",
		16#079c# => X"8326c10d",
		16#079d# => X"13068d00",
		16#079e# => X"13071700",
		16#079f# => X"e3ceb76d",
		16#07a0# => X"83278101",
		16#07a1# => X"2322bd01",
		16#07a2# => X"b38ddd00",
		16#07a3# => X"2320fd00",
		16#07a4# => X"232eb10d",
		16#07a5# => X"232ce10c",
		16#07a6# => X"93067000",
		16#07a7# => X"130d0600",
		16#07a8# => X"63d0e602",
		16#07a9# => X"1306410d",
		16#07aa# => X"93050900",
		16#07ab# => X"13850900",
		16#07ac# => X"ef80906a",
		16#07ad# => X"63040500",
		16#07ae# => X"6f10500c",
		16#07af# => X"130dc10f",
		16#07b0# => X"b38a6a41",
		16#07b1# => X"63505007",
		16#07b2# => X"930d0001",
		16#07b3# => X"13087000",
		16#07b4# => X"83278101",
		16#07b5# => X"0327810d",
		16#07b6# => X"8326c10d",
		16#07b7# => X"2320fd00",
		16#07b8# => X"13071700",
		16#07b9# => X"13068d00",
		16#07ba# => X"e3c05d6d",
		16#07bb# => X"23225d01",
		16#07bc# => X"b38ada00",
		16#07bd# => X"232e510d",
		16#07be# => X"232ce10c",
		16#07bf# => X"93067000",
		16#07c0# => X"130d0600",
		16#07c1# => X"63d0e602",
		16#07c2# => X"1306410d",
		16#07c3# => X"93050900",
		16#07c4# => X"13850900",
		16#07c5# => X"ef805064",
		16#07c6# => X"63040500",
		16#07c7# => X"6f101006",
		16#07c8# => X"130dc10f",
		16#07c9# => X"13770410",
		16#07ca# => X"832dc10d",
		16#07cb# => X"e31e076a",
		16#07cc# => X"8327810d",
		16#07cd# => X"3303bb01",
		16#07ce# => X"23209d00",
		16#07cf# => X"93871700",
		16#07d0# => X"23226d01",
		16#07d1# => X"232e610c",
		16#07d2# => X"232cf10c",
		16#07d3# => X"13077000",
		16#07d4# => X"130d8d00",
		16#07d5# => X"6344f700",
		16#07d6# => X"6f108015",
		16#07d7# => X"1306410d",
		16#07d8# => X"93050900",
		16#07d9# => X"13850900",
		16#07da# => X"ef80105f",
		16#07db# => X"63040500",
		16#07dc# => X"6f10d000",
		16#07dd# => X"130dc10f",
		16#07de# => X"6f108013",
		16#07df# => X"13640401",
		16#07e0# => X"93770402",
		16#07e1# => X"638e0704",
		16#07e2# => X"130c7c00",
		16#07e3# => X"137c8cff",
		16#07e4# => X"93078c00",
		16#07e5# => X"832c0c00",
		16#07e6# => X"032c4c00",
		16#07e7# => X"232ef100",
		16#07e8# => X"635e0c00",
		16#07e9# => X"b30c9041",
		16#07ea# => X"b3379001",
		16#07eb# => X"330c8041",
		16#07ec# => X"330cfc40",
		16#07ed# => X"9307d002",
		16#07ee# => X"a30bf10a",
		16#07ef# => X"9307f0ff",
		16#07f0# => X"e31afb38",
		16#07f1# => X"e31c0c40",
		16#07f2# => X"93079000",
		16#07f3# => X"e3e89741",
		16#07f4# => X"938c0c03",
		16#07f5# => X"a30f9119",
		16#07f6# => X"9304f119",
		16#07f7# => X"6f00903d",
		16#07f8# => X"93074c00",
		16#07f9# => X"232ef100",
		16#07fa# => X"93770401",
		16#07fb# => X"63880700",
		16#07fc# => X"832c0c00",
		16#07fd# => X"13dcfc41",
		16#07fe# => X"6ff09ffa",
		16#07ff# => X"93770404",
		16#0800# => X"832c0c00",
		16#0801# => X"63880700",
		16#0802# => X"939c0c01",
		16#0803# => X"93dc0c41",
		16#0804# => X"6ff05ffe",
		16#0805# => X"93770420",
		16#0806# => X"e38e07fc",
		16#0807# => X"939c8c01",
		16#0808# => X"93dc8c41",
		16#0809# => X"6ff01ffd",
		16#080a# => X"93778400",
		16#080b# => X"638a070a",
		16#080c# => X"93074c00",
		16#080d# => X"232ef100",
		16#080e# => X"83270c00",
		16#080f# => X"03a60700",
		16#0810# => X"83a64700",
		16#0811# => X"03a78700",
		16#0812# => X"83a7c700",
		16#0813# => X"2320c10e",
		16#0814# => X"2322d10e",
		16#0815# => X"2324e10e",
		16#0816# => X"1305010e",
		16#0817# => X"2326f10e",
		16#0818# => X"ef405016",
		16#0819# => X"232ea10a",
		16#081a# => X"93072000",
		16#081b# => X"6310f50c",
		16#081c# => X"8327010e",
		16#081d# => X"93050109",
		16#081e# => X"1305010a",
		16#081f# => X"2320f10a",
		16#0820# => X"8327410e",
		16#0821# => X"23280108",
		16#0822# => X"232a0108",
		16#0823# => X"2322f10a",
		16#0824# => X"8327810e",
		16#0825# => X"232c0108",
		16#0826# => X"232e0108",
		16#0827# => X"2324f10a",
		16#0828# => X"8327c10e",
		16#0829# => X"2326f10a",
		16#082a# => X"efd0c023",
		16#082b# => X"63560500",
		16#082c# => X"9307d002",
		16#082d# => X"a30bf10a",
		16#082e# => X"0327c100",
		16#082f# => X"93077004",
		16#0830# => X"63c0e706",
		16#0831# => X"b7440110",
		16#0832# => X"9384448f",
		16#0833# => X"1374f4f7",
		16#0834# => X"23280100",
		16#0835# => X"130b3000",
		16#0836# => X"930a0000",
		16#0837# => X"6f00902e",
		16#0838# => X"130c7c00",
		16#0839# => X"137c8cff",
		16#083a# => X"83250c00",
		16#083b# => X"03264c00",
		16#083c# => X"93078c00",
		16#083d# => X"1305010a",
		16#083e# => X"232ef100",
		16#083f# => X"eff0d078",
		16#0840# => X"8327010a",
		16#0841# => X"2320f10e",
		16#0842# => X"8327410a",
		16#0843# => X"2322f10e",
		16#0844# => X"8327810a",
		16#0845# => X"2324f10e",
		16#0846# => X"8327c10a",
		16#0847# => X"6ff0dff3",
		16#0848# => X"b7440110",
		16#0849# => X"9384848f",
		16#084a# => X"6ff05ffa",
		16#084b# => X"93071000",
		16#084c# => X"631cf502",
		16#084d# => X"8327c10e",
		16#084e# => X"63d60700",
		16#084f# => X"9307d002",
		16#0850# => X"a30bf10a",
		16#0851# => X"0327c100",
		16#0852# => X"93077004",
		16#0853# => X"63c8e700",
		16#0854# => X"b7440110",
		16#0855# => X"9384c48f",
		16#0856# => X"6ff05ff7",
		16#0857# => X"b7440110",
		16#0858# => X"93840490",
		16#0859# => X"6ff09ff6",
		16#085a# => X"8327c100",
		16#085b# => X"93fbf7fd",
		16#085c# => X"93071004",
		16#085d# => X"6390fb06",
		16#085e# => X"8326c100",
		16#085f# => X"93070003",
		16#0860# => X"230cf10a",
		16#0861# => X"13071006",
		16#0862# => X"93078005",
		16#0863# => X"6394e600",
		16#0864# => X"93078007",
		16#0865# => X"a30cf10a",
		16#0866# => X"93073006",
		16#0867# => X"13642400",
		16#0868# => X"63de6749",
		16#0869# => X"93051b00",
		16#086a# => X"13850900",
		16#086b# => X"ef40d030",
		16#086c# => X"93040500",
		16#086d# => X"631a0548",
		16#086e# => X"8357c900",
		16#086f# => X"93e70704",
		16#0870# => X"2316f900",
		16#0871# => X"8357c900",
		16#0872# => X"93f70704",
		16#0873# => X"638607f6",
		16#0874# => X"6ff08ffb",
		16#0875# => X"9307f0ff",
		16#0876# => X"630cfb46",
		16#0877# => X"93077004",
		16#0878# => X"23280100",
		16#0879# => X"6394fb00",
		16#087a# => X"630a0b46",
		16#087b# => X"032ac10e",
		16#087c# => X"93670410",
		16#087d# => X"2328f102",
		16#087e# => X"23240104",
		16#087f# => X"032e010e",
		16#0880# => X"832d410e",
		16#0881# => X"832c810e",
		16#0882# => X"635a0a00",
		16#0883# => X"b7070080",
		16#0884# => X"33ca4701",
		16#0885# => X"9307d002",
		16#0886# => X"2324f104",
		16#0887# => X"93071004",
		16#0888# => X"6398fb48",
		16#0889# => X"1305010a",
		16#088a# => X"2320c10b",
		16#088b# => X"2324910b",
		16#088c# => X"2322b10b",
		16#088d# => X"2326410b",
		16#088e# => X"ef00010a",
		16#088f# => X"1306c10b",
		16#0890# => X"ef605009",
		16#0891# => X"13860500",
		16#0892# => X"93050500",
		16#0893# => X"1305010a",
		16#0894# => X"eff09063",
		16#0895# => X"8327010a",
		16#0896# => X"13060107",
		16#0897# => X"93050108",
		16#0898# => X"2320f108",
		16#0899# => X"8327410a",
		16#089a# => X"13050109",
		16#089b# => X"23280106",
		16#089c# => X"2322f108",
		16#089d# => X"8327810a",
		16#089e# => X"232a0106",
		16#089f# => X"232c0106",
		16#08a0# => X"2324f108",
		16#08a1# => X"8327c10a",
		16#08a2# => X"2326f108",
		16#08a3# => X"b707fc3f",
		16#08a4# => X"232ef106",
		16#08a5# => X"efd0001b",
		16#08a6# => X"03280109",
		16#08a7# => X"03264109",
		16#08a8# => X"83268109",
		16#08a9# => X"832cc109",
		16#08aa# => X"93050109",
		16#08ab# => X"1305010a",
		16#08ac# => X"2320010b",
		16#08ad# => X"232c0105",
		16#08ae# => X"2322c10a",
		16#08af# => X"232ac104",
		16#08b0# => X"2324d10a",
		16#08b1# => X"2326d104",
		16#08b2# => X"2326910b",
		16#08b3# => X"23280108",
		16#08b4# => X"232a0108",
		16#08b5# => X"232c0108",
		16#08b6# => X"232e0108",
		16#08b7# => X"efc0d05d",
		16#08b8# => X"8326c104",
		16#08b9# => X"03264105",
		16#08ba# => X"03288105",
		16#08bb# => X"63160500",
		16#08bc# => X"13071000",
		16#08bd# => X"232ee10a",
		16#08be# => X"8327c100",
		16#08bf# => X"13071006",
		16#08c0# => X"6394e736",
		16#08c1# => X"374c0110",
		16#08c2# => X"130c4c90",
		16#08c3# => X"130efbff",
		16#08c4# => X"938d0400",
		16#08c5# => X"b7070340",
		16#08c6# => X"93050109",
		16#08c7# => X"232ac108",
		16#08c8# => X"1305010a",
		16#08c9# => X"13060108",
		16#08ca# => X"232cc105",
		16#08cb# => X"23280109",
		16#08cc# => X"2326f108",
		16#08cd# => X"232cd108",
		16#08ce# => X"232e9109",
		16#08cf# => X"23200108",
		16#08d0# => X"23220108",
		16#08d1# => X"23240108",
		16#08d2# => X"efd0c00f",
		16#08d3# => X"0326010a",
		16#08d4# => X"8326410a",
		16#08d5# => X"1305010a",
		16#08d6# => X"232ac104",
		16#08d7# => X"2326d104",
		16#08d8# => X"eff05024",
		16#08d9# => X"93050500",
		16#08da# => X"130a0500",
		16#08db# => X"1305010a",
		16#08dc# => X"832c810a",
		16#08dd# => X"832ac10a",
		16#08de# => X"eff01039",
		16#08df# => X"8327010a",
		16#08e0# => X"03264105",
		16#08e1# => X"8326c104",
		16#08e2# => X"2328f106",
		16#08e3# => X"8327410a",
		16#08e4# => X"2320c108",
		16#08e5# => X"93050108",
		16#08e6# => X"232af106",
		16#08e7# => X"8327810a",
		16#08e8# => X"13060107",
		16#08e9# => X"13050109",
		16#08ea# => X"232cf106",
		16#08eb# => X"8327c10a",
		16#08ec# => X"23249109",
		16#08ed# => X"23265109",
		16#08ee# => X"232ef106",
		16#08ef# => X"2322d108",
		16#08f0# => X"efe0004e",
		16#08f1# => X"b3054c01",
		16#08f2# => X"83c50500",
		16#08f3# => X"032e8105",
		16#08f4# => X"832ac109",
		16#08f5# => X"938d1d00",
		16#08f6# => X"83220109",
		16#08f7# => X"832f4109",
		16#08f8# => X"032f8109",
		16#08f9# => X"2326c105",
		16#08fa# => X"a38fbdfe",
		16#08fb# => X"9307f0ff",
		16#08fc# => X"938c0a00",
		16#08fd# => X"6308fe06",
		16#08fe# => X"130efeff",
		16#08ff# => X"93050109",
		16#0900# => X"1305010a",
		16#0901# => X"2326e107",
		16#0902# => X"2324f107",
		16#0903# => X"23225106",
		16#0904# => X"2320c107",
		16#0905# => X"2320510a",
		16#0906# => X"232e5104",
		16#0907# => X"2322f10b",
		16#0908# => X"232cf105",
		16#0909# => X"2324e10b",
		16#090a# => X"232ae105",
		16#090b# => X"2326510b",
		16#090c# => X"23280108",
		16#090d# => X"232a0108",
		16#090e# => X"232c0108",
		16#090f# => X"232e0108",
		16#0910# => X"efc09047",
		16#0911# => X"83264105",
		16#0912# => X"03268105",
		16#0913# => X"0328c105",
		16#0914# => X"032e0106",
		16#0915# => X"83224106",
		16#0916# => X"832f8106",
		16#0917# => X"032fc106",
		16#0918# => X"e31a05ea",
		16#0919# => X"b70cfe3f",
		16#091a# => X"93050109",
		16#091b# => X"1305010a",
		16#091c# => X"2320510a",
		16#091d# => X"232e5104",
		16#091e# => X"2322f10b",
		16#091f# => X"232cf105",
		16#0920# => X"2324e10b",
		16#0921# => X"232ae105",
		16#0922# => X"2326510b",
		16#0923# => X"23280108",
		16#0924# => X"232a0108",
		16#0925# => X"232c0108",
		16#0926# => X"232e9109",
		16#0927# => X"efc0904e",
		16#0928# => X"6344a004",
		16#0929# => X"8322c105",
		16#092a# => X"832f8105",
		16#092b# => X"032f4105",
		16#092c# => X"93050109",
		16#092d# => X"1305010a",
		16#092e# => X"2320510a",
		16#092f# => X"2322f10b",
		16#0930# => X"2324e10b",
		16#0931# => X"2326510b",
		16#0932# => X"23280108",
		16#0933# => X"232a0108",
		16#0934# => X"232c0108",
		16#0935# => X"232e9109",
		16#0936# => X"efc0103e",
		16#0937# => X"6310051c",
		16#0938# => X"137a1a00",
		16#0939# => X"630c0a1a",
		16#093a# => X"0346fc00",
		16#093b# => X"2326b10d",
		16#093c# => X"93050003",
		16#093d# => X"8326c10c",
		16#093e# => X"9387f6ff",
		16#093f# => X"2326f10c",
		16#0940# => X"83c7f6ff",
		16#0941# => X"6388c716",
		16#0942# => X"13069003",
		16#0943# => X"6398c716",
		16#0944# => X"8347ac00",
		16#0945# => X"a38ff6fe",
		16#0946# => X"138a0d00",
		16#0947# => X"13077004",
		16#0948# => X"330a9a40",
		16#0949# => X"832cc10b",
		16#094a# => X"639aeb2a",
		16#094b# => X"1307d0ff",
		16#094c# => X"63c4ec00",
		16#094d# => X"63589b33",
		16#094e# => X"8327c100",
		16#094f# => X"9387e7ff",
		16#0950# => X"2326f100",
		16#0951# => X"8327c100",
		16#0952# => X"938afcff",
		16#0953# => X"232e510b",
		16#0954# => X"93f6f7fd",
		16#0955# => X"93051004",
		16#0956# => X"0347c100",
		16#0957# => X"13060000",
		16#0958# => X"6398b600",
		16#0959# => X"1307f700",
		16#095a# => X"1377f70f",
		16#095b# => X"13061000",
		16#095c# => X"2302e10c",
		16#095d# => X"9307b002",
		16#095e# => X"63d80a00",
		16#095f# => X"930a1000",
		16#0960# => X"b38a9a41",
		16#0961# => X"9307d002",
		16#0962# => X"a302f10c",
		16#0963# => X"93079000",
		16#0964# => X"63dc5729",
		16#0965# => X"930b310d",
		16#0966# => X"938c0b00",
		16#0967# => X"930d9000",
		16#0968# => X"9305a000",
		16#0969# => X"13850a00",
		16#096a# => X"ef000113",
		16#096b# => X"13050503",
		16#096c# => X"a38fabfe",
		16#096d# => X"9305a000",
		16#096e# => X"13850a00",
		16#096f# => X"ef008109",
		16#0970# => X"138cfbff",
		16#0971# => X"930a0500",
		16#0972# => X"63c2ad24",
		16#0973# => X"930a0503",
		16#0974# => X"938bebff",
		16#0975# => X"a30f5cff",
		16#0976# => X"9307610c",
		16#0977# => X"63ec9b23",
		16#0978# => X"1307410c",
		16#0979# => X"b387e740",
		16#097a# => X"2320f104",
		16#097b# => X"338b4701",
		16#097c# => X"93071000",
		16#097d# => X"63c64701",
		16#097e# => X"93771400",
		16#097f# => X"63860700",
		16#0980# => X"83274102",
		16#0981# => X"330bfb00",
		16#0982# => X"1374f4bf",
		16#0983# => X"93670410",
		16#0984# => X"2328f102",
		16#0985# => X"130c0000",
		16#0986# => X"930b0000",
		16#0987# => X"930c0000",
		16#0988# => X"83278104",
		16#0989# => X"63860700",
		16#098a# => X"1307d002",
		16#098b# => X"a30be10a",
		16#098c# => X"03240103",
		16#098d# => X"930a0000",
		16#098e# => X"6ff00feb",
		16#098f# => X"23280100",
		16#0990# => X"9304c113",
		16#0991# => X"6ff09fba",
		16#0992# => X"2328a100",
		16#0993# => X"6ff01fba",
		16#0994# => X"23280100",
		16#0995# => X"130b6000",
		16#0996# => X"6ff05fb9",
		16#0997# => X"23286101",
		16#0998# => X"130b1000",
		16#0999# => X"6ff09fb8",
		16#099a# => X"374c0110",
		16#099b# => X"130c8c91",
		16#099c# => X"6ff0dfc9",
		16#099d# => X"a38fb6fe",
		16#099e# => X"6ff0dfe7",
		16#099f# => X"93871700",
		16#09a0# => X"93f7f70f",
		16#09a1# => X"6ff01fe9",
		16#09a2# => X"130a1a00",
		16#09a3# => X"a30feafe",
		16#09a4# => X"b3874a41",
		16#09a5# => X"e3da07fe",
		16#09a6# => X"6ff05fe8",
		16#09a7# => X"8327c104",
		16#09a8# => X"138a0d00",
		16#09a9# => X"13070003",
		16#09aa# => X"b38afd00",
		16#09ab# => X"6ff05ffe",
		16#09ac# => X"93076004",
		16#09ad# => X"638efb00",
		16#09ae# => X"93075004",
		16#09af# => X"930a1b00",
		16#09b0# => X"6384fb00",
		16#09b1# => X"930a0b00",
		16#09b2# => X"13062000",
		16#09b3# => X"6f00c000",
		16#09b4# => X"930a0b00",
		16#09b5# => X"13063000",
		16#09b6# => X"9307010c",
		16#09b7# => X"1308c10c",
		16#09b8# => X"1307c10b",
		16#09b9# => X"93860a00",
		16#09ba# => X"9305010a",
		16#09bb# => X"13850900",
		16#09bc# => X"2320c10b",
		16#09bd# => X"2326c105",
		16#09be# => X"2322b10b",
		16#09bf# => X"2324910b",
		16#09c0# => X"2326410b",
		16#09c1# => X"ef30c066",
		16#09c2# => X"93077004",
		16#09c3# => X"93040500",
		16#09c4# => X"032ec104",
		16#09c5# => X"6396fb00",
		16#09c6# => X"93771400",
		16#09c7# => X"6380070a",
		16#09c8# => X"93076004",
		16#09c9# => X"338c5401",
		16#09ca# => X"639efb04",
		16#09cb# => X"03c70400",
		16#09cc# => X"93070003",
		16#09cd# => X"6314f704",
		16#09ce# => X"93050109",
		16#09cf# => X"1305010a",
		16#09d0# => X"2320c10b",
		16#09d1# => X"2326c105",
		16#09d2# => X"2322b10b",
		16#09d3# => X"2324910b",
		16#09d4# => X"2326410b",
		16#09d5# => X"23280108",
		16#09d6# => X"232a0108",
		16#09d7# => X"232c0108",
		16#09d8# => X"232e0108",
		16#09d9# => X"efc05015",
		16#09da# => X"032ec104",
		16#09db# => X"63080500",
		16#09dc# => X"93071000",
		16#09dd# => X"b38a5741",
		16#09de# => X"232e510b",
		16#09df# => X"8327c10b",
		16#09e0# => X"330cfc00",
		16#09e1# => X"93050109",
		16#09e2# => X"1305010a",
		16#09e3# => X"2320c10b",
		16#09e4# => X"2322b10b",
		16#09e5# => X"2324910b",
		16#09e6# => X"2326410b",
		16#09e7# => X"23280108",
		16#09e8# => X"232a0108",
		16#09e9# => X"232c0108",
		16#09ea# => X"232e0108",
		16#09eb# => X"efc0d010",
		16#09ec# => X"13070003",
		16#09ed# => X"631e0500",
		16#09ee# => X"2326810d",
		16#09ef# => X"032ac10c",
		16#09f0# => X"6ff0dfd5",
		16#09f1# => X"93861700",
		16#09f2# => X"2326d10c",
		16#09f3# => X"2380e700",
		16#09f4# => X"8327c10c",
		16#09f5# => X"e3e887ff",
		16#09f6# => X"6ff05ffe",
		16#09f7# => X"13076004",
		16#09f8# => X"e392ebd6",
		16#09f9# => X"63549007",
		16#09fa# => X"63160b00",
		16#09fb# => X"13771400",
		16#09fc# => X"6306070c",
		16#09fd# => X"83274102",
		16#09fe# => X"3387fc00",
		16#09ff# => X"330beb00",
		16#0a00# => X"93076006",
		16#0a01# => X"2326f100",
		16#0a02# => X"6f008009",
		16#0a03# => X"930b0c00",
		16#0a04# => X"6ff01fd9",
		16#0a05# => X"938b1b00",
		16#0a06# => X"03c7fbff",
		16#0a07# => X"93871700",
		16#0a08# => X"a38fe7fe",
		16#0a09# => X"6ff09fdb",
		16#0a0a# => X"1307610c",
		16#0a0b# => X"63180600",
		16#0a0c# => X"93070003",
		16#0a0d# => X"2303f10c",
		16#0a0e# => X"1307710c",
		16#0a0f# => X"938a0a03",
		16#0a10# => X"93071700",
		16#0a11# => X"23005701",
		16#0a12# => X"6ff09fd9",
		16#0a13# => X"63160b00",
		16#0a14# => X"13771400",
		16#0a15# => X"63080706",
		16#0a16# => X"83274102",
		16#0a17# => X"13871700",
		16#0a18# => X"6ff0dff9",
		16#0a19# => X"63c04c03",
		16#0a1a# => X"13771400",
		16#0a1b# => X"138b0c00",
		16#0a1c# => X"63060700",
		16#0a1d# => X"83274102",
		16#0a1e# => X"338bfc00",
		16#0a1f# => X"93077006",
		16#0a20# => X"6ff05ff8",
		16#0a21# => X"83274102",
		16#0a22# => X"330bfa00",
		16#0a23# => X"93077006",
		16#0a24# => X"2326f100",
		16#0a25# => X"63469001",
		16#0a26# => X"33039b41",
		16#0a27# => X"130b1300",
		16#0a28# => X"937b0440",
		16#0a29# => X"130c0000",
		16#0a2a# => X"e38c0bd6",
		16#0a2b# => X"930b0000",
		16#0a2c# => X"e35890d7",
		16#0a2d# => X"9306f00f",
		16#0a2e# => X"6f00c003",
		16#0a2f# => X"138b0c00",
		16#0a30# => X"6ff01ff4",
		16#0a31# => X"93076006",
		16#0a32# => X"2326f100",
		16#0a33# => X"130b1000",
		16#0a34# => X"6ff01ffd",
		16#0a35# => X"63569703",
		16#0a36# => X"83274101",
		16#0a37# => X"b38cec40",
		16#0a38# => X"03c71700",
		16#0a39# => X"63080702",
		16#0a3a# => X"93871700",
		16#0a3b# => X"938b1b00",
		16#0a3c# => X"232af100",
		16#0a3d# => X"83274101",
		16#0a3e# => X"03c70700",
		16#0a3f# => X"e31cd7fc",
		16#0a40# => X"83254103",
		16#0a41# => X"33858b01",
		16#0a42# => X"eff09052",
		16#0a43# => X"330b6501",
		16#0a44# => X"6ff01fd1",
		16#0a45# => X"130c1c00",
		16#0a46# => X"6ff0dffd",
		16#0a47# => X"13074c00",
		16#0a48# => X"232ee100",
		16#0a49# => X"13770402",
		16#0a4a# => X"83270c00",
		16#0a4b# => X"63000702",
		16#0a4c# => X"03278102",
		16#0a4d# => X"23a0e700",
		16#0a4e# => X"1357f741",
		16#0a4f# => X"23a2e700",
		16#0a50# => X"032cc101",
		16#0a51# => X"83240102",
		16#0a52# => X"6ff04f89",
		16#0a53# => X"13770401",
		16#0a54# => X"63080700",
		16#0a55# => X"03278102",
		16#0a56# => X"23a0e700",
		16#0a57# => X"6ff05ffe",
		16#0a58# => X"13770404",
		16#0a59# => X"63080700",
		16#0a5a# => X"03578102",
		16#0a5b# => X"2390e700",
		16#0a5c# => X"6ff01ffd",
		16#0a5d# => X"13740420",
		16#0a5e# => X"e30e04fc",
		16#0a5f# => X"03478102",
		16#0a60# => X"2380e700",
		16#0a61# => X"6ff0dffb",
		16#0a62# => X"13640401",
		16#0a63# => X"93770402",
		16#0a64# => X"63880704",
		16#0a65# => X"130c7c00",
		16#0a66# => X"137c8cff",
		16#0a67# => X"93078c00",
		16#0a68# => X"832c0c00",
		16#0a69# => X"032c4c00",
		16#0a6a# => X"232ef100",
		16#0a6b# => X"1374f4bf",
		16#0a6c# => X"93070000",
		16#0a6d# => X"a30b010a",
		16#0a6e# => X"1307f0ff",
		16#0a6f# => X"6302eb1a",
		16#0a70# => X"13070400",
		16#0a71# => X"b3e68c01",
		16#0a72# => X"1374f4f7",
		16#0a73# => X"639a0618",
		16#0a74# => X"630c0b2e",
		16#0a75# => X"13071000",
		16#0a76# => X"6398e718",
		16#0a77# => X"6ff04fdf",
		16#0a78# => X"93074c00",
		16#0a79# => X"232ef100",
		16#0a7a# => X"93770401",
		16#0a7b# => X"63860700",
		16#0a7c# => X"832c0c00",
		16#0a7d# => X"6f000001",
		16#0a7e# => X"93770404",
		16#0a7f# => X"63880700",
		16#0a80# => X"835c0c00",
		16#0a81# => X"130c0000",
		16#0a82# => X"6ff05ffa",
		16#0a83# => X"93770420",
		16#0a84# => X"e38007fe",
		16#0a85# => X"834c0c00",
		16#0a86# => X"6ff0dffe",
		16#0a87# => X"93074c00",
		16#0a88# => X"232ef100",
		16#0a89# => X"b787ffff",
		16#0a8a# => X"93c70783",
		16#0a8b# => X"231cf10a",
		16#0a8c# => X"b7470110",
		16#0a8d# => X"93874790",
		16#0a8e# => X"13078007",
		16#0a8f# => X"832c0c00",
		16#0a90# => X"2322f104",
		16#0a91# => X"130c0000",
		16#0a92# => X"13642400",
		16#0a93# => X"93072000",
		16#0a94# => X"2326e100",
		16#0a95# => X"6ff01ff6",
		16#0a96# => X"93074c00",
		16#0a97# => X"232ef100",
		16#0a98# => X"a30b010a",
		16#0a99# => X"9307f0ff",
		16#0a9a# => X"83240c00",
		16#0a9b# => X"6304fb02",
		16#0a9c# => X"13060b00",
		16#0a9d# => X"93050000",
		16#0a9e# => X"13850400",
		16#0a9f# => X"ef401010",
		16#0aa0# => X"2328a100",
		16#0aa1# => X"630a05e4",
		16#0aa2# => X"330b9540",
		16#0aa3# => X"23280100",
		16#0aa4# => X"6ff08fe4",
		16#0aa5# => X"13850400",
		16#0aa6# => X"efe0dfd7",
		16#0aa7# => X"130b0500",
		16#0aa8# => X"6ff0dffe",
		16#0aa9# => X"13640401",
		16#0aaa# => X"93770402",
		16#0aab# => X"63820702",
		16#0aac# => X"130c7c00",
		16#0aad# => X"137c8cff",
		16#0aae# => X"93078c00",
		16#0aaf# => X"832c0c00",
		16#0ab0# => X"032c4c00",
		16#0ab1# => X"232ef100",
		16#0ab2# => X"93071000",
		16#0ab3# => X"6ff09fee",
		16#0ab4# => X"93074c00",
		16#0ab5# => X"232ef100",
		16#0ab6# => X"93770401",
		16#0ab7# => X"63860700",
		16#0ab8# => X"832c0c00",
		16#0ab9# => X"6f000001",
		16#0aba# => X"93770404",
		16#0abb# => X"63880700",
		16#0abc# => X"835c0c00",
		16#0abd# => X"130c0000",
		16#0abe# => X"6ff01ffd",
		16#0abf# => X"93770420",
		16#0ac0# => X"e38007fe",
		16#0ac1# => X"834c0c00",
		16#0ac2# => X"6ff0dffe",
		16#0ac3# => X"b7470110",
		16#0ac4# => X"93874790",
		16#0ac5# => X"6fe0dffa",
		16#0ac6# => X"93074c00",
		16#0ac7# => X"232ef100",
		16#0ac8# => X"93770401",
		16#0ac9# => X"63860700",
		16#0aca# => X"832c0c00",
		16#0acb# => X"6f000001",
		16#0acc# => X"93770404",
		16#0acd# => X"63880700",
		16#0ace# => X"835c0c00",
		16#0acf# => X"130c0000",
		16#0ad0# => X"6fe09ffa",
		16#0ad1# => X"93770420",
		16#0ad2# => X"e38007fe",
		16#0ad3# => X"834c0c00",
		16#0ad4# => X"6ff0dffe",
		16#0ad5# => X"13070400",
		16#0ad6# => X"93071000",
		16#0ad7# => X"6ff09fe6",
		16#0ad8# => X"13071000",
		16#0ad9# => X"6380e7c6",
		16#0ada# => X"13072000",
		16#0adb# => X"6382e712",
		16#0adc# => X"9307011a",
		16#0add# => X"9316dc01",
		16#0ade# => X"13f77c00",
		16#0adf# => X"93dc3c00",
		16#0ae0# => X"13070703",
		16#0ae1# => X"b3ec9601",
		16#0ae2# => X"135c3c00",
		16#0ae3# => X"a38fe7fe",
		16#0ae4# => X"b3e68c01",
		16#0ae5# => X"9384f7ff",
		16#0ae6# => X"639e0602",
		16#0ae7# => X"93761400",
		16#0ae8# => X"638a0600",
		16#0ae9# => X"93060003",
		16#0aea# => X"6306d700",
		16#0aeb# => X"a38fd4fe",
		16#0aec# => X"9384e7ff",
		16#0aed# => X"9307011a",
		16#0aee# => X"930a0b00",
		16#0aef# => X"23280100",
		16#0af0# => X"338b9740",
		16#0af1# => X"130c0000",
		16#0af2# => X"930b0000",
		16#0af3# => X"930c0000",
		16#0af4# => X"6ff08f91",
		16#0af5# => X"93870400",
		16#0af6# => X"6ff0dff9",
		16#0af7# => X"130a0000",
		16#0af8# => X"930d011a",
		16#0af9# => X"937a0440",
		16#0afa# => X"930b9000",
		16#0afb# => X"1306a000",
		16#0afc# => X"93060000",
		16#0afd# => X"13850c00",
		16#0afe# => X"93050c00",
		16#0aff# => X"efb0400c",
		16#0b00# => X"13050503",
		16#0b01# => X"a38fadfe",
		16#0b02# => X"9384fdff",
		16#0b03# => X"130a1a00",
		16#0b04# => X"638a0a04",
		16#0b05# => X"83274101",
		16#0b06# => X"83c70700",
		16#0b07# => X"6314fa04",
		16#0b08# => X"9307f00f",
		16#0b09# => X"6300fa04",
		16#0b0a# => X"63140c00",
		16#0b0b# => X"63fc9b03",
		16#0b0c# => X"83274103",
		16#0b0d# => X"8325c103",
		16#0b0e# => X"130a0000",
		16#0b0f# => X"b384f440",
		16#0b10# => X"13860700",
		16#0b11# => X"13850400",
		16#0b12# => X"ef608016",
		16#0b13# => X"83274101",
		16#0b14# => X"83c71700",
		16#0b15# => X"63880700",
		16#0b16# => X"83274101",
		16#0b17# => X"93871700",
		16#0b18# => X"232af100",
		16#0b19# => X"13850c00",
		16#0b1a# => X"93050c00",
		16#0b1b# => X"1306a000",
		16#0b1c# => X"93060000",
		16#0b1d# => X"efa01027",
		16#0b1e# => X"138c0500",
		16#0b1f# => X"b3e5a500",
		16#0b20# => X"930c0500",
		16#0b21# => X"e38805f2",
		16#0b22# => X"938d0400",
		16#0b23# => X"6ff01ff6",
		16#0b24# => X"9304011a",
		16#0b25# => X"03274104",
		16#0b26# => X"93f7fc00",
		16#0b27# => X"9384f4ff",
		16#0b28# => X"b307f700",
		16#0b29# => X"83c70700",
		16#0b2a# => X"93dc4c00",
		16#0b2b# => X"2380f400",
		16#0b2c# => X"9317cc01",
		16#0b2d# => X"b3ec9701",
		16#0b2e# => X"135c4c00",
		16#0b2f# => X"b3e78c01",
		16#0b30# => X"e39a07fc",
		16#0b31# => X"6ff01fef",
		16#0b32# => X"9304011a",
		16#0b33# => X"e39407ee",
		16#0b34# => X"13771700",
		16#0b35# => X"e30007ee",
		16#0b36# => X"93070003",
		16#0b37# => X"a30ff118",
		16#0b38# => X"6ff08faf",
		16#0b39# => X"8327c100",
		16#0b3a# => X"e38c072e",
		16#0b3b# => X"8347c100",
		16#0b3c# => X"a30b010a",
		16#0b3d# => X"232e8101",
		16#0b3e# => X"230ef112",
		16#0b3f# => X"6fe01ffd",
		16#0b40# => X"13060601",
		16#0b41# => X"2322dd01",
		16#0b42# => X"232ec10c",
		16#0b43# => X"232cd10c",
		16#0b44# => X"635edf02",
		16#0b45# => X"1306410d",
		16#0b46# => X"93050900",
		16#0b47# => X"13850900",
		16#0b48# => X"232ee105",
		16#0b49# => X"232cc105",
		16#0b4a# => X"232ad105",
		16#0b4b# => X"2326e104",
		16#0b4c# => X"ef808002",
		16#0b4d# => X"e3140524",
		16#0b4e# => X"032fc105",
		16#0b4f# => X"032e8105",
		16#0b50# => X"832e4105",
		16#0b51# => X"0327c104",
		16#0b52# => X"9305c10f",
		16#0b53# => X"130707ff",
		16#0b54# => X"138d0500",
		16#0b55# => X"6fe05fff",
		16#0b56# => X"83258101",
		16#0b57# => X"93860601",
		16#0b58# => X"2322fd00",
		16#0b59# => X"2320bd00",
		16#0b5a# => X"232ed10c",
		16#0b5b# => X"232ce10c",
		16#0b5c# => X"6356ee02",
		16#0b5d# => X"1306410d",
		16#0b5e# => X"93050900",
		16#0b5f# => X"13850900",
		16#0b60# => X"2326c105",
		16#0b61# => X"2324f104",
		16#0b62# => X"ef70107d",
		16#0b63# => X"e318051e",
		16#0b64# => X"032ec104",
		16#0b65# => X"83278104",
		16#0b66# => X"1306c10f",
		16#0b67# => X"938d0dff",
		16#0b68# => X"130d0600",
		16#0b69# => X"6ff08f8c",
		16#0b6a# => X"93860601",
		16#0b6b# => X"2322bd01",
		16#0b6c# => X"232ed10c",
		16#0b6d# => X"232ce10c",
		16#0b6e# => X"6352e802",
		16#0b6f# => X"1306410d",
		16#0b70# => X"93050900",
		16#0b71# => X"13850900",
		16#0b72# => X"23240105",
		16#0b73# => X"ef70d078",
		16#0b74# => X"e316051a",
		16#0b75# => X"03288104",
		16#0b76# => X"1306c10f",
		16#0b77# => X"938a0aff",
		16#0b78# => X"130d0600",
		16#0b79# => X"6ff0cf8e",
		16#0b7a# => X"8327c100",
		16#0b7b# => X"13075006",
		16#0b7c# => X"6354f772",
		16#0b7d# => X"0327010e",
		16#0b7e# => X"93050109",
		16#0b7f# => X"1305010a",
		16#0b80# => X"2320e10a",
		16#0b81# => X"0327410e",
		16#0b82# => X"23280108",
		16#0b83# => X"232a0108",
		16#0b84# => X"2322e10a",
		16#0b85# => X"0327810e",
		16#0b86# => X"232c0108",
		16#0b87# => X"232e0108",
		16#0b88# => X"2324e10a",
		16#0b89# => X"0327c10e",
		16#0b8a# => X"2326e10a",
		16#0b8b# => X"efc0c028",
		16#0b8c# => X"631a0512",
		16#0b8d# => X"b7470110",
		16#0b8e# => X"9387c792",
		16#0b8f# => X"2320fd00",
		16#0b90# => X"93071000",
		16#0b91# => X"2322fd00",
		16#0b92# => X"8327810d",
		16#0b93# => X"938d1d00",
		16#0b94# => X"232eb10d",
		16#0b95# => X"93871700",
		16#0b96# => X"232cf10c",
		16#0b97# => X"13077000",
		16#0b98# => X"130d8d00",
		16#0b99# => X"635ef700",
		16#0b9a# => X"1306410d",
		16#0b9b# => X"93050900",
		16#0b9c# => X"13850900",
		16#0b9d# => X"ef70506e",
		16#0b9e# => X"e3120510",
		16#0b9f# => X"130dc10f",
		16#0ba0# => X"8327c10b",
		16#0ba1# => X"63c64701",
		16#0ba2# => X"93771400",
		16#0ba3# => X"63820722",
		16#0ba4# => X"83278103",
		16#0ba5# => X"03274102",
		16#0ba6# => X"130d8d00",
		16#0ba7# => X"232cfdfe",
		16#0ba8# => X"83274102",
		16#0ba9# => X"232efdfe",
		16#0baa# => X"8327c10d",
		16#0bab# => X"b387e700",
		16#0bac# => X"232ef10c",
		16#0bad# => X"8327810d",
		16#0bae# => X"13077000",
		16#0baf# => X"93871700",
		16#0bb0# => X"232cf10c",
		16#0bb1# => X"635ef700",
		16#0bb2# => X"1306410d",
		16#0bb3# => X"93050900",
		16#0bb4# => X"13850900",
		16#0bb5# => X"ef705068",
		16#0bb6# => X"e312050a",
		16#0bb7# => X"130dc10f",
		16#0bb8# => X"9304faff",
		16#0bb9# => X"6356901c",
		16#0bba# => X"930a0001",
		16#0bbb# => X"930b7000",
		16#0bbc# => X"03268101",
		16#0bbd# => X"8327810d",
		16#0bbe# => X"0327c10d",
		16#0bbf# => X"2320cd00",
		16#0bc0# => X"93871700",
		16#0bc1# => X"93068d00",
		16#0bc2# => X"63c29a02",
		16#0bc3# => X"23229d00",
		16#0bc4# => X"b384e400",
		16#0bc5# => X"232e910c",
		16#0bc6# => X"232cf10c",
		16#0bc7# => X"13077000",
		16#0bc8# => X"138d0600",
		16#0bc9# => X"6356f718",
		16#0bca# => X"6ff04f83",
		16#0bcb# => X"13070701",
		16#0bcc# => X"23225d01",
		16#0bcd# => X"232ee10c",
		16#0bce# => X"232cf10c",
		16#0bcf# => X"63defb00",
		16#0bd0# => X"1306410d",
		16#0bd1# => X"93050900",
		16#0bd2# => X"13850900",
		16#0bd3# => X"ef70d060",
		16#0bd4# => X"e3160502",
		16#0bd5# => X"9306c10f",
		16#0bd6# => X"938404ff",
		16#0bd7# => X"138d0600",
		16#0bd8# => X"6ff01ff9",
		16#0bd9# => X"0327c10b",
		16#0bda# => X"634ae01c",
		16#0bdb# => X"b7470110",
		16#0bdc# => X"9387c792",
		16#0bdd# => X"2320fd00",
		16#0bde# => X"93071000",
		16#0bdf# => X"2322fd00",
		16#0be0# => X"8327810d",
		16#0be1# => X"938d1d00",
		16#0be2# => X"232eb10d",
		16#0be3# => X"93871700",
		16#0be4# => X"232cf10c",
		16#0be5# => X"13077000",
		16#0be6# => X"130d8d00",
		16#0be7# => X"635ef700",
		16#0be8# => X"1306410d",
		16#0be9# => X"93050900",
		16#0bea# => X"13850900",
		16#0beb# => X"ef70d05a",
		16#0bec# => X"6316057c",
		16#0bed# => X"130dc10f",
		16#0bee# => X"8327c10b",
		16#0bef# => X"63980700",
		16#0bf0# => X"63160a00",
		16#0bf1# => X"93771400",
		16#0bf2# => X"6384070e",
		16#0bf3# => X"83278103",
		16#0bf4# => X"03274102",
		16#0bf5# => X"93088d00",
		16#0bf6# => X"2320fd00",
		16#0bf7# => X"83274102",
		16#0bf8# => X"2322fd00",
		16#0bf9# => X"8327c10d",
		16#0bfa# => X"b387e700",
		16#0bfb# => X"232ef10c",
		16#0bfc# => X"8327810d",
		16#0bfd# => X"13077000",
		16#0bfe# => X"93871700",
		16#0bff# => X"232cf10c",
		16#0c00# => X"635ef700",
		16#0c01# => X"1306410d",
		16#0c02# => X"93050900",
		16#0c03# => X"13850900",
		16#0c04# => X"ef709054",
		16#0c05# => X"63140576",
		16#0c06# => X"9308c10f",
		16#0c07# => X"832ac10b",
		16#0c08# => X"63d00a06",
		16#0c09# => X"b30a5041",
		16#0c0a# => X"13870800",
		16#0c0b# => X"930b0001",
		16#0c0c# => X"130c7000",
		16#0c0d# => X"03268101",
		16#0c0e# => X"8327810d",
		16#0c0f# => X"8326c10d",
		16#0c10# => X"2320c700",
		16#0c11# => X"93871700",
		16#0c12# => X"93888800",
		16#0c13# => X"63cc5b0b",
		16#0c14# => X"23225701",
		16#0c15# => X"b38ada00",
		16#0c16# => X"232e510d",
		16#0c17# => X"232cf10c",
		16#0c18# => X"13077000",
		16#0c19# => X"635ef700",
		16#0c1a# => X"1306410d",
		16#0c1b# => X"93050900",
		16#0c1c# => X"13850900",
		16#0c1d# => X"ef70504e",
		16#0c1e# => X"63120570",
		16#0c1f# => X"9308c10f",
		16#0c20# => X"8327c10d",
		16#0c21# => X"23a09800",
		16#0c22# => X"23a24801",
		16#0c23# => X"b3874701",
		16#0c24# => X"232ef10c",
		16#0c25# => X"8327810d",
		16#0c26# => X"13077000",
		16#0c27# => X"138d8800",
		16#0c28# => X"93871700",
		16#0c29# => X"232cf10c",
		16#0c2a# => X"6354f700",
		16#0c2b# => X"6fe01feb",
		16#0c2c# => X"13744400",
		16#0c2d# => X"63140466",
		16#0c2e# => X"032dc102",
		16#0c2f# => X"83270103",
		16#0c30# => X"6354fd00",
		16#0c31# => X"138d0700",
		16#0c32# => X"83278102",
		16#0c33# => X"b387a701",
		16#0c34# => X"2324f102",
		16#0c35# => X"8327c10d",
		16#0c36# => X"638c0700",
		16#0c37# => X"1306410d",
		16#0c38# => X"93050900",
		16#0c39# => X"13850900",
		16#0c3a# => X"ef701047",
		16#0c3b# => X"63180568",
		16#0c3c# => X"83270101",
		16#0c3d# => X"232c010c",
		16#0c3e# => X"639c076c",
		16#0c3f# => X"130dc10f",
		16#0c40# => X"6ff01f84",
		16#0c41# => X"93860601",
		16#0c42# => X"23227701",
		16#0c43# => X"232ed10c",
		16#0c44# => X"232cf10c",
		16#0c45# => X"635efc00",
		16#0c46# => X"1306410d",
		16#0c47# => X"93050900",
		16#0c48# => X"13850900",
		16#0c49# => X"ef705043",
		16#0c4a# => X"631a0564",
		16#0c4b# => X"9308c10f",
		16#0c4c# => X"938a0aff",
		16#0c4d# => X"13870800",
		16#0c4e# => X"6ff0dfef",
		16#0c4f# => X"938a0c00",
		16#0c50# => X"63549a01",
		16#0c51# => X"930a0a00",
		16#0c52# => X"63525005",
		16#0c53# => X"0327810d",
		16#0c54# => X"b38dba01",
		16#0c55# => X"23209d00",
		16#0c56# => X"13071700",
		16#0c57# => X"23225d01",
		16#0c58# => X"232eb10d",
		16#0c59# => X"232ce10c",
		16#0c5a# => X"93067000",
		16#0c5b# => X"130d8d00",
		16#0c5c# => X"63dee600",
		16#0c5d# => X"1306410d",
		16#0c5e# => X"93050900",
		16#0c5f# => X"13850900",
		16#0c60# => X"ef70903d",
		16#0c61# => X"631c055e",
		16#0c62# => X"130dc10f",
		16#0c63# => X"63d40a00",
		16#0c64# => X"930a0000",
		16#0c65# => X"b38a5c41",
		16#0c66# => X"635e5005",
		16#0c67# => X"130b0001",
		16#0c68# => X"930d7000",
		16#0c69# => X"83278101",
		16#0c6a# => X"0327810d",
		16#0c6b# => X"8326c10d",
		16#0c6c# => X"2320fd00",
		16#0c6d# => X"13071700",
		16#0c6e# => X"13068d00",
		16#0c6f# => X"634c5b19",
		16#0c70# => X"23225d01",
		16#0c71# => X"b38ada00",
		16#0c72# => X"232e510d",
		16#0c73# => X"232ce10c",
		16#0c74# => X"93067000",
		16#0c75# => X"130d0600",
		16#0c76# => X"63dee600",
		16#0c77# => X"1306410d",
		16#0c78# => X"93050900",
		16#0c79# => X"13850900",
		16#0c7a# => X"ef701037",
		16#0c7b# => X"63180558",
		16#0c7c# => X"130dc10f",
		16#0c7d# => X"93770440",
		16#0c7e# => X"b38a9401",
		16#0c7f# => X"63800702",
		16#0c80# => X"130b7000",
		16#0c81# => X"b38d4401",
		16#0c82# => X"63920b18",
		16#0c83# => X"63120c18",
		16#0c84# => X"b3874401",
		16#0c85# => X"63f45701",
		16#0c86# => X"938a0700",
		16#0c87# => X"8327c10b",
		16#0c88# => X"63c64701",
		16#0c89# => X"93771400",
		16#0c8a# => X"638a0704",
		16#0c8b# => X"83278103",
		16#0c8c# => X"03274102",
		16#0c8d# => X"130d8d00",
		16#0c8e# => X"232cfdfe",
		16#0c8f# => X"83274102",
		16#0c90# => X"232efdfe",
		16#0c91# => X"8327c10d",
		16#0c92# => X"b387e700",
		16#0c93# => X"232ef10c",
		16#0c94# => X"8327810d",
		16#0c95# => X"13077000",
		16#0c96# => X"93871700",
		16#0c97# => X"232cf10c",
		16#0c98# => X"635ef700",
		16#0c99# => X"1306410d",
		16#0c9a# => X"93050900",
		16#0c9b# => X"13850900",
		16#0c9c# => X"ef70902e",
		16#0c9d# => X"63140550",
		16#0c9e# => X"130dc10f",
		16#0c9f# => X"b3844401",
		16#0ca0# => X"b3875441",
		16#0ca1# => X"8324c10b",
		16#0ca2# => X"b3049a40",
		16#0ca3# => X"63d49700",
		16#0ca4# => X"93840700",
		16#0ca5# => X"63549004",
		16#0ca6# => X"8327c10d",
		16#0ca7# => X"23205d01",
		16#0ca8# => X"23229d00",
		16#0ca9# => X"b387f400",
		16#0caa# => X"232ef10c",
		16#0cab# => X"8327810d",
		16#0cac# => X"13077000",
		16#0cad# => X"130d8d00",
		16#0cae# => X"93871700",
		16#0caf# => X"232cf10c",
		16#0cb0# => X"635ef700",
		16#0cb1# => X"1306410d",
		16#0cb2# => X"93050900",
		16#0cb3# => X"13850900",
		16#0cb4# => X"ef709028",
		16#0cb5# => X"6314054a",
		16#0cb6# => X"130dc10f",
		16#0cb7# => X"93870400",
		16#0cb8# => X"63d40400",
		16#0cb9# => X"93070000",
		16#0cba# => X"8324c10b",
		16#0cbb# => X"b3049a40",
		16#0cbc# => X"b384f440",
		16#0cbd# => X"e35e90da",
		16#0cbe# => X"930a0001",
		16#0cbf# => X"930b7000",
		16#0cc0# => X"03268101",
		16#0cc1# => X"8327810d",
		16#0cc2# => X"0327c10d",
		16#0cc3# => X"2320cd00",
		16#0cc4# => X"93871700",
		16#0cc5# => X"93068d00",
		16#0cc6# => X"e3da9abe",
		16#0cc7# => X"13070701",
		16#0cc8# => X"23225d01",
		16#0cc9# => X"232ee10c",
		16#0cca# => X"232cf10c",
		16#0ccb# => X"63defb00",
		16#0ccc# => X"1306410d",
		16#0ccd# => X"93050900",
		16#0cce# => X"13850900",
		16#0ccf# => X"ef70d021",
		16#0cd0# => X"631e0542",
		16#0cd1# => X"9306c10f",
		16#0cd2# => X"938404ff",
		16#0cd3# => X"138d0600",
		16#0cd4# => X"6ff01ffb",
		16#0cd5# => X"93860601",
		16#0cd6# => X"23226d01",
		16#0cd7# => X"232ed10c",
		16#0cd8# => X"232ce10c",
		16#0cd9# => X"63deed00",
		16#0cda# => X"1306410d",
		16#0cdb# => X"93050900",
		16#0cdc# => X"13850900",
		16#0cdd# => X"ef70501e",
		16#0cde# => X"63120540",
		16#0cdf# => X"1306c10f",
		16#0ce0# => X"938a0aff",
		16#0ce1# => X"130d0600",
		16#0ce2# => X"6ff0dfe1",
		16#0ce3# => X"63020c0e",
		16#0ce4# => X"130cfcff",
		16#0ce5# => X"8327c103",
		16#0ce6# => X"03274103",
		16#0ce7# => X"130d8d00",
		16#0ce8# => X"232cfdfe",
		16#0ce9# => X"83274103",
		16#0cea# => X"232efdfe",
		16#0ceb# => X"8327c10d",
		16#0cec# => X"b387e700",
		16#0ced# => X"232ef10c",
		16#0cee# => X"8327810d",
		16#0cef# => X"93871700",
		16#0cf0# => X"232cf10c",
		16#0cf1# => X"635efb00",
		16#0cf2# => X"1306410d",
		16#0cf3# => X"93050900",
		16#0cf4# => X"13850900",
		16#0cf5# => X"ef705018",
		16#0cf6# => X"6312053a",
		16#0cf7# => X"130dc10f",
		16#0cf8# => X"83274101",
		16#0cf9# => X"33875d41",
		16#0cfa# => X"83c70700",
		16#0cfb# => X"6354f700",
		16#0cfc# => X"93070700",
		16#0cfd# => X"6356f004",
		16#0cfe# => X"0327c10d",
		16#0cff# => X"23205d01",
		16#0d00# => X"2322fd00",
		16#0d01# => X"3387e700",
		16#0d02# => X"232ee10c",
		16#0d03# => X"0327810d",
		16#0d04# => X"130d8d00",
		16#0d05# => X"13071700",
		16#0d06# => X"232ce10c",
		16#0d07# => X"6352eb02",
		16#0d08# => X"1306410d",
		16#0d09# => X"93050900",
		16#0d0a# => X"13850900",
		16#0d0b# => X"2326f100",
		16#0d0c# => X"ef709012",
		16#0d0d# => X"63140534",
		16#0d0e# => X"8327c100",
		16#0d0f# => X"130dc10f",
		16#0d10# => X"13870700",
		16#0d11# => X"63d40700",
		16#0d12# => X"13070000",
		16#0d13# => X"83274101",
		16#0d14# => X"13080001",
		16#0d15# => X"83c70700",
		16#0d16# => X"b387e740",
		16#0d17# => X"6346f006",
		16#0d18# => X"83274101",
		16#0d19# => X"83c70700",
		16#0d1a# => X"b38afa00",
		16#0d1b# => X"6ff0dfd9",
		16#0d1c# => X"83274101",
		16#0d1d# => X"938bfbff",
		16#0d1e# => X"9387f7ff",
		16#0d1f# => X"232af100",
		16#0d20# => X"6ff05ff1",
		16#0d21# => X"93860601",
		16#0d22# => X"23220d01",
		16#0d23# => X"232ed10c",
		16#0d24# => X"232ce10c",
		16#0d25# => X"6356eb02",
		16#0d26# => X"1306410d",
		16#0d27# => X"93050900",
		16#0d28# => X"13850900",
		16#0d29# => X"23240105",
		16#0d2a# => X"2326f100",
		16#0d2b# => X"ef70d00a",
		16#0d2c# => X"6316052c",
		16#0d2d# => X"03288104",
		16#0d2e# => X"8327c100",
		16#0d2f# => X"1306c10f",
		16#0d30# => X"938707ff",
		16#0d31# => X"130d0600",
		16#0d32# => X"83258101",
		16#0d33# => X"0327810d",
		16#0d34# => X"8326c10d",
		16#0d35# => X"2320bd00",
		16#0d36# => X"13071700",
		16#0d37# => X"13068d00",
		16#0d38# => X"e342f8fa",
		16#0d39# => X"2322fd00",
		16#0d3a# => X"b387d700",
		16#0d3b# => X"232ef10c",
		16#0d3c# => X"232ce10c",
		16#0d3d# => X"130d0600",
		16#0d3e# => X"e354ebf6",
		16#0d3f# => X"1306410d",
		16#0d40# => X"93050900",
		16#0d41# => X"13850900",
		16#0d42# => X"ef701005",
		16#0d43# => X"63180526",
		16#0d44# => X"130dc10f",
		16#0d45# => X"6ff0dff4",
		16#0d46# => X"8327810d",
		16#0d47# => X"13071000",
		16#0d48# => X"23209d00",
		16#0d49# => X"938d1d00",
		16#0d4a# => X"93871700",
		16#0d4b# => X"930b8d00",
		16#0d4c# => X"63464701",
		16#0d4d# => X"93761400",
		16#0d4e# => X"6386061c",
		16#0d4f# => X"13071000",
		16#0d50# => X"2322ed00",
		16#0d51# => X"232eb10d",
		16#0d52# => X"232cf10c",
		16#0d53# => X"13077000",
		16#0d54# => X"635ef700",
		16#0d55# => X"1306410d",
		16#0d56# => X"93050900",
		16#0d57# => X"13850900",
		16#0d58# => X"ef70807f",
		16#0d59# => X"631c0520",
		16#0d5a# => X"930bc10f",
		16#0d5b# => X"83278103",
		16#0d5c# => X"03274102",
		16#0d5d# => X"938b8b00",
		16#0d5e# => X"23acfbfe",
		16#0d5f# => X"83274102",
		16#0d60# => X"23aefbfe",
		16#0d61# => X"8327c10d",
		16#0d62# => X"b387e700",
		16#0d63# => X"232ef10c",
		16#0d64# => X"8327810d",
		16#0d65# => X"13077000",
		16#0d66# => X"93871700",
		16#0d67# => X"232cf10c",
		16#0d68# => X"635ef700",
		16#0d69# => X"1306410d",
		16#0d6a# => X"93050900",
		16#0d6b# => X"13850900",
		16#0d6c# => X"ef70807a",
		16#0d6d# => X"6314051c",
		16#0d6e# => X"930bc10f",
		16#0d6f# => X"8327010e",
		16#0d70# => X"93050109",
		16#0d71# => X"1305010a",
		16#0d72# => X"2320f10a",
		16#0d73# => X"8327410e",
		16#0d74# => X"930afaff",
		16#0d75# => X"23280108",
		16#0d76# => X"2322f10a",
		16#0d77# => X"8327810e",
		16#0d78# => X"232a0108",
		16#0d79# => X"232c0108",
		16#0d7a# => X"2324f10a",
		16#0d7b# => X"8327c10e",
		16#0d7c# => X"232e0108",
		16#0d7d# => X"2326f10a",
		16#0d7e# => X"efb0102c",
		16#0d7f# => X"63060508",
		16#0d80# => X"8327c10d",
		16#0d81# => X"0327810d",
		16#0d82# => X"93841400",
		16#0d83# => X"9387f7ff",
		16#0d84# => X"b3874701",
		16#0d85# => X"13071700",
		16#0d86# => X"23a09b00",
		16#0d87# => X"23a25b01",
		16#0d88# => X"232ef10c",
		16#0d89# => X"232ce10c",
		16#0d8a# => X"93077000",
		16#0d8b# => X"938b8b00",
		16#0d8c# => X"63dee700",
		16#0d8d# => X"1306410d",
		16#0d8e# => X"93050900",
		16#0d8f# => X"13850900",
		16#0d90# => X"ef708071",
		16#0d91# => X"631c0512",
		16#0d92# => X"930bc10f",
		16#0d93# => X"9307410c",
		16#0d94# => X"23a0fb00",
		16#0d95# => X"83270104",
		16#0d96# => X"03270104",
		16#0d97# => X"138d8b00",
		16#0d98# => X"23a2fb00",
		16#0d99# => X"8327c10d",
		16#0d9a# => X"b387e700",
		16#0d9b# => X"232ef10c",
		16#0d9c# => X"8327810d",
		16#0d9d# => X"13077000",
		16#0d9e# => X"93871700",
		16#0d9f# => X"232cf10c",
		16#0da0# => X"e358f7a2",
		16#0da1# => X"6fe09f8d",
		16#0da2# => X"e35250fd",
		16#0da3# => X"93040001",
		16#0da4# => X"130c7000",
		16#0da5# => X"03268101",
		16#0da6# => X"0327810d",
		16#0da7# => X"8327c10d",
		16#0da8# => X"23a0cb00",
		16#0da9# => X"13071700",
		16#0daa# => X"93868b00",
		16#0dab# => X"63c05403",
		16#0dac# => X"b387fa00",
		16#0dad# => X"23a25b01",
		16#0dae# => X"232ef10c",
		16#0daf# => X"232ce10c",
		16#0db0# => X"93077000",
		16#0db1# => X"938b0600",
		16#0db2# => X"6ff09ff6",
		16#0db3# => X"93870701",
		16#0db4# => X"23a29b00",
		16#0db5# => X"232ef10c",
		16#0db6# => X"232ce10c",
		16#0db7# => X"635eec00",
		16#0db8# => X"1306410d",
		16#0db9# => X"93050900",
		16#0dba# => X"13850900",
		16#0dbb# => X"ef70c066",
		16#0dbc# => X"63160508",
		16#0dbd# => X"9306c10f",
		16#0dbe# => X"938a0aff",
		16#0dbf# => X"938b0600",
		16#0dc0# => X"6ff05ff9",
		16#0dc1# => X"2322ed00",
		16#0dc2# => X"232eb10d",
		16#0dc3# => X"232cf10c",
		16#0dc4# => X"13077000",
		16#0dc5# => X"e35cf7f2",
		16#0dc6# => X"6ff0dff1",
		16#0dc7# => X"8327c102",
		16#0dc8# => X"03270103",
		16#0dc9# => X"3384e740",
		16#0dca# => X"e3588098",
		16#0dcb# => X"b7440110",
		16#0dcc# => X"930a0001",
		16#0dcd# => X"938444cc",
		16#0dce# => X"930b7000",
		16#0dcf# => X"8327810d",
		16#0dd0# => X"23209d00",
		16#0dd1# => X"0327c10d",
		16#0dd2# => X"93871700",
		16#0dd3# => X"63c68a04",
		16#0dd4# => X"23228d00",
		16#0dd5# => X"3304e400",
		16#0dd6# => X"232e810c",
		16#0dd7# => X"232cf10c",
		16#0dd8# => X"13077000",
		16#0dd9# => X"e35af794",
		16#0dda# => X"1306410d",
		16#0ddb# => X"93050900",
		16#0ddc# => X"13850900",
		16#0ddd# => X"ef70405e",
		16#0dde# => X"e3000594",
		16#0ddf# => X"83270101",
		16#0de0# => X"63940700",
		16#0de1# => X"6fe01fa4",
		16#0de2# => X"93850700",
		16#0de3# => X"13850900",
		16#0de4# => X"ef00d020",
		16#0de5# => X"6fe01fa3",
		16#0de6# => X"13070701",
		16#0de7# => X"23225d01",
		16#0de8# => X"232ee10c",
		16#0de9# => X"232cf10c",
		16#0dea# => X"130d8d00",
		16#0deb# => X"63defb00",
		16#0dec# => X"1306410d",
		16#0ded# => X"93050900",
		16#0dee# => X"13850900",
		16#0def# => X"ef70c059",
		16#0df0# => X"e31e05fa",
		16#0df1# => X"130dc10f",
		16#0df2# => X"130404ff",
		16#0df3# => X"6ff01ff7",
		16#0df4# => X"83250101",
		16#0df5# => X"13850900",
		16#0df6# => X"ef00501c",
		16#0df7# => X"6ff01f92",
		16#0df8# => X"8327c10d",
		16#0df9# => X"63940700",
		16#0dfa# => X"6fe0df9d",
		16#0dfb# => X"1306410d",
		16#0dfc# => X"93050900",
		16#0dfd# => X"13850900",
		16#0dfe# => X"ef700056",
		16#0dff# => X"6fe09f9c",
		16#0e00# => X"93060600",
		16#0e01# => X"13860500",
		16#0e02# => X"93050500",
		16#0e03# => X"03a5c181",
		16#0e04# => X"6fe04f83",
		16#0e05# => X"83d7c500",
		16#0e06# => X"130101b8",
		16#0e07# => X"232c8146",
		16#0e08# => X"93f7d7ff",
		16#0e09# => X"231af100",
		16#0e0a# => X"83a74506",
		16#0e0b# => X"13840500",
		16#0e0c# => X"232a9146",
		16#0e0d# => X"2326f106",
		16#0e0e# => X"83d7e500",
		16#0e0f# => X"23282147",
		16#0e10# => X"232e1146",
		16#0e11# => X"231bf100",
		16#0e12# => X"83a7c501",
		16#0e13# => X"13090500",
		16#0e14# => X"23200102",
		16#0e15# => X"2322f102",
		16#0e16# => X"83a74502",
		16#0e17# => X"93058100",
		16#0e18# => X"2326f102",
		16#0e19# => X"93070107",
		16#0e1a# => X"2324f100",
		16#0e1b# => X"232cf100",
		16#0e1c# => X"93070040",
		16#0e1d# => X"2328f100",
		16#0e1e# => X"232ef100",
		16#0e1f# => X"efd09ffc",
		16#0e20# => X"93040500",
		16#0e21# => X"634c0500",
		16#0e22# => X"93058100",
		16#0e23# => X"13050900",
		16#0e24# => X"ef00c04b",
		16#0e25# => X"63040500",
		16#0e26# => X"9304f0ff",
		16#0e27# => X"83574101",
		16#0e28# => X"93f70704",
		16#0e29# => X"63880700",
		16#0e2a# => X"8357c400",
		16#0e2b# => X"93e70704",
		16#0e2c# => X"2316f400",
		16#0e2d# => X"8320c147",
		16#0e2e# => X"03248147",
		16#0e2f# => X"13850400",
		16#0e30# => X"03290147",
		16#0e31# => X"83244147",
		16#0e32# => X"13010148",
		16#0e33# => X"67800000",
		16#0e34# => X"130101fe",
		16#0e35# => X"232c8100",
		16#0e36# => X"232a9100",
		16#0e37# => X"23282101",
		16#0e38# => X"232e1100",
		16#0e39# => X"23263101",
		16#0e3a# => X"13090500",
		16#0e3b# => X"93840500",
		16#0e3c# => X"13040600",
		16#0e3d# => X"63080500",
		16#0e3e# => X"83278503",
		16#0e3f# => X"63940700",
		16#0e40# => X"ef00805e",
		16#0e41# => X"83278401",
		16#0e42# => X"2324f400",
		16#0e43# => X"8357c400",
		16#0e44# => X"93f78700",
		16#0e45# => X"638a0708",
		16#0e46# => X"83270401",
		16#0e47# => X"63860708",
		16#0e48# => X"8317c400",
		16#0e49# => X"93f9f40f",
		16#0e4a# => X"93f4f40f",
		16#0e4b# => X"13972701",
		16#0e4c# => X"6356070a",
		16#0e4d# => X"83270401",
		16#0e4e# => X"03250400",
		16#0e4f# => X"3305f540",
		16#0e50# => X"83274401",
		16#0e51# => X"634af500",
		16#0e52# => X"93050400",
		16#0e53# => X"13050900",
		16#0e54# => X"ef00c03f",
		16#0e55# => X"63120506",
		16#0e56# => X"83278400",
		16#0e57# => X"13051500",
		16#0e58# => X"9387f7ff",
		16#0e59# => X"2324f400",
		16#0e5a# => X"83270400",
		16#0e5b# => X"13871700",
		16#0e5c# => X"2320e400",
		16#0e5d# => X"23803701",
		16#0e5e# => X"83274401",
		16#0e5f# => X"638ca700",
		16#0e60# => X"8357c400",
		16#0e61# => X"93f71700",
		16#0e62# => X"638a0702",
		16#0e63# => X"9307a000",
		16#0e64# => X"6396f402",
		16#0e65# => X"93050400",
		16#0e66# => X"13050900",
		16#0e67# => X"ef00003b",
		16#0e68# => X"630e0500",
		16#0e69# => X"6f004001",
		16#0e6a# => X"93050400",
		16#0e6b# => X"13050900",
		16#0e6c# => X"ef000006",
		16#0e6d# => X"e30605f6",
		16#0e6e# => X"9304f0ff",
		16#0e6f# => X"8320c101",
		16#0e70# => X"03248101",
		16#0e71# => X"13850400",
		16#0e72# => X"03290101",
		16#0e73# => X"83244101",
		16#0e74# => X"8329c100",
		16#0e75# => X"13010102",
		16#0e76# => X"67800000",
		16#0e77# => X"37270000",
		16#0e78# => X"b3e7e700",
		16#0e79# => X"2316f400",
		16#0e7a# => X"83274406",
		16#0e7b# => X"37e7ffff",
		16#0e7c# => X"1307f7ff",
		16#0e7d# => X"b3f7e700",
		16#0e7e# => X"2322f406",
		16#0e7f# => X"6ff09ff3",
		16#0e80# => X"13860500",
		16#0e81# => X"93050500",
		16#0e82# => X"03a5c181",
		16#0e83# => X"6ff05fec",
		16#0e84# => X"130101ff",
		16#0e85# => X"23229100",
		16#0e86# => X"93040500",
		16#0e87# => X"03a5c181",
		16#0e88# => X"23248100",
		16#0e89# => X"23261100",
		16#0e8a# => X"13840500",
		16#0e8b# => X"63080500",
		16#0e8c# => X"83278503",
		16#0e8d# => X"63940700",
		16#0e8e# => X"ef00004b",
		16#0e8f# => X"0317c400",
		16#0e90# => X"93170701",
		16#0e91# => X"93d70701",
		16#0e92# => X"93f68700",
		16#0e93# => X"639e0606",
		16#0e94# => X"93f60701",
		16#0e95# => X"63960602",
		16#0e96# => X"93079000",
		16#0e97# => X"23a0f400",
		16#0e98# => X"13670704",
		16#0e99# => X"2316e400",
		16#0e9a# => X"1305f0ff",
		16#0e9b# => X"8320c100",
		16#0e9c# => X"03248100",
		16#0e9d# => X"83244100",
		16#0e9e# => X"13010101",
		16#0e9f# => X"67800000",
		16#0ea0# => X"93f74700",
		16#0ea1# => X"638c0702",
		16#0ea2# => X"83250403",
		16#0ea3# => X"638c0500",
		16#0ea4# => X"93070404",
		16#0ea5# => X"6386f500",
		16#0ea6# => X"13850400",
		16#0ea7# => X"ef000070",
		16#0ea8# => X"23280402",
		16#0ea9# => X"8357c400",
		16#0eaa# => X"23220400",
		16#0eab# => X"93f7b7fd",
		16#0eac# => X"2316f400",
		16#0ead# => X"83270401",
		16#0eae# => X"2320f400",
		16#0eaf# => X"8357c400",
		16#0eb0# => X"93e78700",
		16#0eb1# => X"2316f400",
		16#0eb2# => X"83270401",
		16#0eb3# => X"63900702",
		16#0eb4# => X"8357c400",
		16#0eb5# => X"13070020",
		16#0eb6# => X"93f70728",
		16#0eb7# => X"6388e700",
		16#0eb8# => X"93050400",
		16#0eb9# => X"13850400",
		16#0eba# => X"ef30000e",
		16#0ebb# => X"8357c400",
		16#0ebc# => X"13f71700",
		16#0ebd# => X"630c0702",
		16#0ebe# => X"83274401",
		16#0ebf# => X"23240400",
		16#0ec0# => X"b307f040",
		16#0ec1# => X"232cf400",
		16#0ec2# => X"83270401",
		16#0ec3# => X"13050000",
		16#0ec4# => X"e39e07f4",
		16#0ec5# => X"8317c400",
		16#0ec6# => X"13f70708",
		16#0ec7# => X"e30807f4",
		16#0ec8# => X"93e70704",
		16#0ec9# => X"2316f400",
		16#0eca# => X"6ff01ff4",
		16#0ecb# => X"93f72700",
		16#0ecc# => X"13070000",
		16#0ecd# => X"63940700",
		16#0ece# => X"03274401",
		16#0ecf# => X"2324e400",
		16#0ed0# => X"6ff09ffc",
		16#0ed1# => X"8397c500",
		16#0ed2# => X"130101fe",
		16#0ed3# => X"232c8100",
		16#0ed4# => X"13970701",
		16#0ed5# => X"13570701",
		16#0ed6# => X"232a9100",
		16#0ed7# => X"232e1100",
		16#0ed8# => X"23282101",
		16#0ed9# => X"23263101",
		16#0eda# => X"93768700",
		16#0edb# => X"93040500",
		16#0edc# => X"13840500",
		16#0edd# => X"639c0616",
		16#0ede# => X"37170000",
		16#0edf# => X"13070780",
		16#0ee0# => X"b3e7e700",
		16#0ee1# => X"03a74500",
		16#0ee2# => X"2396f500",
		16#0ee3# => X"6346e002",
		16#0ee4# => X"03a7c503",
		16#0ee5# => X"6342e002",
		16#0ee6# => X"13050000",
		16#0ee7# => X"8320c101",
		16#0ee8# => X"03248101",
		16#0ee9# => X"83244101",
		16#0eea# => X"03290101",
		16#0eeb# => X"8329c100",
		16#0eec# => X"13010102",
		16#0eed# => X"67800000",
		16#0eee# => X"03278402",
		16#0eef# => X"e30e07fc",
		16#0ef0# => X"03a90400",
		16#0ef1# => X"93963701",
		16#0ef2# => X"23a00400",
		16#0ef3# => X"8325c401",
		16#0ef4# => X"63d8060c",
		16#0ef5# => X"03260405",
		16#0ef6# => X"8357c400",
		16#0ef7# => X"93f74700",
		16#0ef8# => X"638e0700",
		16#0ef9# => X"83274400",
		16#0efa# => X"3306f640",
		16#0efb# => X"83270403",
		16#0efc# => X"63860700",
		16#0efd# => X"8327c403",
		16#0efe# => X"3306f640",
		16#0eff# => X"83278402",
		16#0f00# => X"8325c401",
		16#0f01# => X"93060000",
		16#0f02# => X"13850400",
		16#0f03# => X"e7800700",
		16#0f04# => X"9307f0ff",
		16#0f05# => X"8356c400",
		16#0f06# => X"6312f502",
		16#0f07# => X"83a70400",
		16#0f08# => X"1307d001",
		16#0f09# => X"636cf70a",
		16#0f0a# => X"37074020",
		16#0f0b# => X"13071700",
		16#0f0c# => X"3357f700",
		16#0f0d# => X"13771700",
		16#0f0e# => X"6302070a",
		16#0f0f# => X"b7f7ffff",
		16#0f10# => X"9387f77f",
		16#0f11# => X"03270401",
		16#0f12# => X"b3f7d700",
		16#0f13# => X"93970701",
		16#0f14# => X"93d70741",
		16#0f15# => X"2320e400",
		16#0f16# => X"2316f400",
		16#0f17# => X"23220400",
		16#0f18# => X"13973701",
		16#0f19# => X"635c0700",
		16#0f1a# => X"9307f0ff",
		16#0f1b# => X"6316f500",
		16#0f1c# => X"83a70400",
		16#0f1d# => X"63940700",
		16#0f1e# => X"2328a404",
		16#0f1f# => X"83250403",
		16#0f20# => X"23a02401",
		16#0f21# => X"e38a05f0",
		16#0f22# => X"93070404",
		16#0f23# => X"6386f500",
		16#0f24# => X"13850400",
		16#0f25# => X"ef008050",
		16#0f26# => X"23280402",
		16#0f27# => X"6ff0dfef",
		16#0f28# => X"13060000",
		16#0f29# => X"93061000",
		16#0f2a# => X"13850400",
		16#0f2b# => X"e7000700",
		16#0f2c# => X"9307f0ff",
		16#0f2d# => X"13060500",
		16#0f2e# => X"e310f5f2",
		16#0f2f# => X"83a70400",
		16#0f30# => X"e38c07f0",
		16#0f31# => X"1307d001",
		16#0f32# => X"6386e700",
		16#0f33# => X"13076001",
		16#0f34# => X"6392e706",
		16#0f35# => X"23a02401",
		16#0f36# => X"6ff01fec",
		16#0f37# => X"93e70604",
		16#0f38# => X"2316f400",
		16#0f39# => X"1305f0ff",
		16#0f3a# => X"6ff05feb",
		16#0f3b# => X"83a90501",
		16#0f3c# => X"e38409ea",
		16#0f3d# => X"03a90500",
		16#0f3e# => X"13773700",
		16#0f3f# => X"23a03501",
		16#0f40# => X"33093941",
		16#0f41# => X"93070000",
		16#0f42# => X"63140700",
		16#0f43# => X"83a74501",
		16#0f44# => X"2324f400",
		16#0f45# => X"e35220e9",
		16#0f46# => X"83274402",
		16#0f47# => X"8325c401",
		16#0f48# => X"93060900",
		16#0f49# => X"13860900",
		16#0f4a# => X"13850400",
		16#0f4b# => X"e7800700",
		16#0f4c# => X"6348a000",
		16#0f4d# => X"8357c400",
		16#0f4e# => X"93e70704",
		16#0f4f# => X"6ff05ffa",
		16#0f50# => X"b389a900",
		16#0f51# => X"3309a940",
		16#0f52# => X"6ff0dffc",
		16#0f53# => X"130101fe",
		16#0f54# => X"232c8100",
		16#0f55# => X"232e1100",
		16#0f56# => X"13040500",
		16#0f57# => X"630c0500",
		16#0f58# => X"83278503",
		16#0f59# => X"63980700",
		16#0f5a# => X"2326b100",
		16#0f5b# => X"ef00c017",
		16#0f5c# => X"8325c100",
		16#0f5d# => X"8397c500",
		16#0f5e# => X"638c0700",
		16#0f5f# => X"13050400",
		16#0f60# => X"03248101",
		16#0f61# => X"8320c101",
		16#0f62# => X"13010102",
		16#0f63# => X"6ff09fdb",
		16#0f64# => X"8320c101",
		16#0f65# => X"03248101",
		16#0f66# => X"13050000",
		16#0f67# => X"13010102",
		16#0f68# => X"67800000",
		16#0f69# => X"93050500",
		16#0f6a# => X"631a0500",
		16#0f6b# => X"03a58181",
		16#0f6c# => X"b7450010",
		16#0f6d# => X"9385c5d4",
		16#0f6e# => X"6f005034",
		16#0f6f# => X"03a5c181",
		16#0f70# => X"6ff0dff8",
		16#0f71# => X"13050000",
		16#0f72# => X"67800000",
		16#0f73# => X"b7c50010",
		16#0f74# => X"938545d3",
		16#0f75# => X"6f009032",
		16#0f76# => X"130101ff",
		16#0f77# => X"23248100",
		16#0f78# => X"23261100",
		16#0f79# => X"13040500",
		16#0f7a# => X"2316b500",
		16#0f7b# => X"2317c500",
		16#0f7c# => X"23200500",
		16#0f7d# => X"23220500",
		16#0f7e# => X"23240500",
		16#0f7f# => X"23220506",
		16#0f80# => X"23280500",
		16#0f81# => X"232a0500",
		16#0f82# => X"232c0500",
		16#0f83# => X"13068000",
		16#0f84# => X"93050000",
		16#0f85# => X"1305c505",
		16#0f86# => X"ef30406c",
		16#0f87# => X"b7970010",
		16#0f88# => X"938787c5",
		16#0f89# => X"2320f402",
		16#0f8a# => X"b7970010",
		16#0f8b# => X"938707cb",
		16#0f8c# => X"2322f402",
		16#0f8d# => X"b7970010",
		16#0f8e# => X"938747d3",
		16#0f8f# => X"2324f402",
		16#0f90# => X"b7970010",
		16#0f91# => X"9387c7d8",
		16#0f92# => X"232e8400",
		16#0f93# => X"2326f402",
		16#0f94# => X"8320c100",
		16#0f95# => X"03248100",
		16#0f96# => X"13010101",
		16#0f97# => X"67800000",
		16#0f98# => X"13050000",
		16#0f99# => X"67800000",
		16#0f9a# => X"130101ff",
		16#0f9b# => X"23202101",
		16#0f9c# => X"13890500",
		16#0f9d# => X"23248100",
		16#0f9e# => X"93058006",
		16#0f9f# => X"13040500",
		16#0fa0# => X"1305f9ff",
		16#0fa1# => X"23261100",
		16#0fa2# => X"23229100",
		16#0fa3# => X"efe0407a",
		16#0fa4# => X"93054507",
		16#0fa5# => X"93040500",
		16#0fa6# => X"13050400",
		16#0fa7# => X"ef20d061",
		16#0fa8# => X"13040500",
		16#0fa9# => X"63000502",
		16#0faa# => X"23200500",
		16#0fab# => X"23222501",
		16#0fac# => X"1305c500",
		16#0fad# => X"2324a400",
		16#0fae# => X"13868406",
		16#0faf# => X"93050000",
		16#0fb0# => X"ef30c061",
		16#0fb1# => X"13050400",
		16#0fb2# => X"8320c100",
		16#0fb3# => X"03248100",
		16#0fb4# => X"83244100",
		16#0fb5# => X"03290100",
		16#0fb6# => X"13010101",
		16#0fb7# => X"67800000",
		16#0fb8# => X"03a58181",
		16#0fb9# => X"6ff09fee",
		16#0fba# => X"83278503",
		16#0fbb# => X"639e0706",
		16#0fbc# => X"130101ff",
		16#0fbd# => X"b7470010",
		16#0fbe# => X"23261100",
		16#0fbf# => X"23248100",
		16#0fc0# => X"9387c7dc",
		16#0fc1# => X"232ef502",
		16#0fc2# => X"93073000",
		16#0fc3# => X"2322f52e",
		16#0fc4# => X"9307c52e",
		16#0fc5# => X"13040500",
		16#0fc6# => X"2324f52e",
		16#0fc7# => X"2320052e",
		16#0fc8# => X"03254500",
		16#0fc9# => X"13060000",
		16#0fca# => X"93054000",
		16#0fcb# => X"eff0dfea",
		16#0fcc# => X"03258400",
		16#0fcd# => X"13061000",
		16#0fce# => X"93059000",
		16#0fcf# => X"eff0dfe9",
		16#0fd0# => X"0325c400",
		16#0fd1# => X"13062000",
		16#0fd2# => X"93052001",
		16#0fd3# => X"eff0dfe8",
		16#0fd4# => X"93071000",
		16#0fd5# => X"232cf402",
		16#0fd6# => X"8320c100",
		16#0fd7# => X"03248100",
		16#0fd8# => X"13010101",
		16#0fd9# => X"67800000",
		16#0fda# => X"67800000",
		16#0fdb# => X"130101ff",
		16#0fdc# => X"23229100",
		16#0fdd# => X"83a48181",
		16#0fde# => X"23202101",
		16#0fdf# => X"23261100",
		16#0fe0# => X"83a78403",
		16#0fe1# => X"23248100",
		16#0fe2# => X"13090500",
		16#0fe3# => X"63960700",
		16#0fe4# => X"13850400",
		16#0fe5# => X"eff05ff5",
		16#0fe6# => X"9384042e",
		16#0fe7# => X"03a48400",
		16#0fe8# => X"83a74400",
		16#0fe9# => X"9387f7ff",
		16#0fea# => X"63da0700",
		16#0feb# => X"83a70400",
		16#0fec# => X"638e0700",
		16#0fed# => X"83a40400",
		16#0fee# => X"6ff05ffe",
		16#0fef# => X"0317c400",
		16#0ff0# => X"63040704",
		16#0ff1# => X"13048406",
		16#0ff2# => X"6ff0dffd",
		16#0ff3# => X"93054000",
		16#0ff4# => X"13050900",
		16#0ff5# => X"eff05fe9",
		16#0ff6# => X"23a0a400",
		16#0ff7# => X"e31c05fc",
		16#0ff8# => X"9307c000",
		16#0ff9# => X"2320f900",
		16#0ffa# => X"13040000",
		16#0ffb# => X"13050400",
		16#0ffc# => X"8320c100",
		16#0ffd# => X"03248100",
		16#0ffe# => X"83244100",
		16#0fff# => X"03290100",
		16#1000# => X"13010101",
		16#1001# => X"67800000",
		16#1002# => X"b707ffff",
		16#1003# => X"93871700",
		16#1004# => X"23220406",
		16#1005# => X"23200400",
		16#1006# => X"23220400",
		16#1007# => X"23240400",
		16#1008# => X"2326f400",
		16#1009# => X"23280400",
		16#100a# => X"232a0400",
		16#100b# => X"232c0400",
		16#100c# => X"13068000",
		16#100d# => X"93050000",
		16#100e# => X"1305c405",
		16#100f# => X"ef30004a",
		16#1010# => X"23280402",
		16#1011# => X"232a0402",
		16#1012# => X"23220404",
		16#1013# => X"23240404",
		16#1014# => X"6ff0dff9",
		16#1015# => X"67800000",
		16#1016# => X"67800000",
		16#1017# => X"67800000",
		16#1018# => X"67800000",
		16#1019# => X"03a5c181",
		16#101a# => X"b7450010",
		16#101b# => X"938545dc",
		16#101c# => X"6f00c07e",
		16#101d# => X"03a5c181",
		16#101e# => X"b7450010",
		16#101f# => X"938505e6",
		16#1020# => X"6f00c07d",
		16#1021# => X"130101fd",
		16#1022# => X"23202103",
		16#1023# => X"37590110",
		16#1024# => X"23248102",
		16#1025# => X"23229102",
		16#1026# => X"232e3101",
		16#1027# => X"2326b100",
		16#1028# => X"23261102",
		16#1029# => X"93090500",
		16#102a# => X"1309c9e0",
		16#102b# => X"ef30c050",
		16#102c# => X"83278900",
		16#102d# => X"8325c100",
		16#102e# => X"83a44700",
		16#102f# => X"b7170000",
		16#1030# => X"1384f7fe",
		16#1031# => X"93f4c4ff",
		16#1032# => X"3304b440",
		16#1033# => X"33049400",
		16#1034# => X"1354c400",
		16#1035# => X"1304f4ff",
		16#1036# => X"1314c400",
		16#1037# => X"6356f402",
		16#1038# => X"13850900",
		16#1039# => X"ef30804d",
		16#103a# => X"13050000",
		16#103b# => X"8320c102",
		16#103c# => X"03248102",
		16#103d# => X"83244102",
		16#103e# => X"03290102",
		16#103f# => X"8329c101",
		16#1040# => X"13010103",
		16#1041# => X"67800000",
		16#1042# => X"93050000",
		16#1043# => X"13850900",
		16#1044# => X"ef409017",
		16#1045# => X"83278900",
		16#1046# => X"b3879700",
		16#1047# => X"e312f5fc",
		16#1048# => X"b3058040",
		16#1049# => X"13850900",
		16#104a# => X"ef401016",
		16#104b# => X"9307f0ff",
		16#104c# => X"631ef502",
		16#104d# => X"93050000",
		16#104e# => X"13850900",
		16#104f# => X"ef40d014",
		16#1050# => X"03278900",
		16#1051# => X"9306f000",
		16#1052# => X"b307e540",
		16#1053# => X"e3daf6f8",
		16#1054# => X"83a60182",
		16#1055# => X"93e71700",
		16#1056# => X"2322f700",
		16#1057# => X"3305d540",
		16#1058# => X"b7560110",
		16#1059# => X"23a4a626",
		16#105a# => X"6ff09ff7",
		16#105b# => X"83278900",
		16#105c# => X"b3848440",
		16#105d# => X"37570110",
		16#105e# => X"93e41400",
		16#105f# => X"23a29700",
		16#1060# => X"83278726",
		16#1061# => X"13850900",
		16#1062# => X"33848740",
		16#1063# => X"23248726",
		16#1064# => X"ef30c042",
		16#1065# => X"13051000",
		16#1066# => X"6ff05ff5",
		16#1067# => X"638c0524",
		16#1068# => X"130101ff",
		16#1069# => X"23248100",
		16#106a# => X"23229100",
		16#106b# => X"13040500",
		16#106c# => X"93840500",
		16#106d# => X"23261100",
		16#106e# => X"ef300040",
		16#106f# => X"03a5c4ff",
		16#1070# => X"37560110",
		16#1071# => X"938684ff",
		16#1072# => X"9377e5ff",
		16#1073# => X"1308c6e0",
		16#1074# => X"b385f600",
		16#1075# => X"03a74500",
		16#1076# => X"03288800",
		16#1077# => X"1306c6e0",
		16#1078# => X"1377c7ff",
		16#1079# => X"13751500",
		16#107a# => X"6310b806",
		16#107b# => X"b387e700",
		16#107c# => X"63100502",
		16#107d# => X"03a784ff",
		16#107e# => X"b386e640",
		16#107f# => X"83a58600",
		16#1080# => X"b387e700",
		16#1081# => X"03a7c600",
		16#1082# => X"23a6e500",
		16#1083# => X"2324b700",
		16#1084# => X"13e71700",
		16#1085# => X"23a2e600",
		16#1086# => X"03a74182",
		16#1087# => X"2324d600",
		16#1088# => X"63e8e700",
		16#1089# => X"83a54184",
		16#108a# => X"13050400",
		16#108b# => X"eff09fe5",
		16#108c# => X"13050400",
		16#108d# => X"03248100",
		16#108e# => X"8320c100",
		16#108f# => X"83244100",
		16#1090# => X"13010101",
		16#1091# => X"6f308037",
		16#1092# => X"23a2e500",
		16#1093# => X"13080000",
		16#1094# => X"63160502",
		16#1095# => X"03a584ff",
		16#1096# => X"b7580110",
		16#1097# => X"938848e1",
		16#1098# => X"b386a640",
		16#1099# => X"b387a700",
		16#109a# => X"03a58600",
		16#109b# => X"6306150b",
		16#109c# => X"83a8c600",
		16#109d# => X"23261501",
		16#109e# => X"23a4a800",
		16#109f# => X"3385e500",
		16#10a0# => X"03254500",
		16#10a1# => X"13751500",
		16#10a2# => X"63180502",
		16#10a3# => X"b387e700",
		16#10a4# => X"03a78500",
		16#10a5# => X"63160808",
		16#10a6# => X"37550110",
		16#10a7# => X"130545e1",
		16#10a8# => X"6310a708",
		16#10a9# => X"232ad600",
		16#10aa# => X"2328d600",
		16#10ab# => X"23a6e600",
		16#10ac# => X"23a4e600",
		16#10ad# => X"13081000",
		16#10ae# => X"13e71700",
		16#10af# => X"23a2e600",
		16#10b0# => X"3387f600",
		16#10b1# => X"2320f700",
		16#10b2# => X"e31408f6",
		16#10b3# => X"1307f01f",
		16#10b4# => X"6360f706",
		16#10b5# => X"93d73700",
		16#10b6# => X"93d52740",
		16#10b7# => X"13071000",
		16#10b8# => X"3317b700",
		16#10b9# => X"83254600",
		16#10ba# => X"93871700",
		16#10bb# => X"93973700",
		16#10bc# => X"b307f600",
		16#10bd# => X"3367b700",
		16#10be# => X"2322e600",
		16#10bf# => X"03a70700",
		16#10c0# => X"138687ff",
		16#10c1# => X"23a6c600",
		16#10c2# => X"23a4e600",
		16#10c3# => X"23a0d700",
		16#10c4# => X"2326d700",
		16#10c5# => X"6ff0dff1",
		16#10c6# => X"13081000",
		16#10c7# => X"6ff01ff6",
		16#10c8# => X"83a5c500",
		16#10c9# => X"2326b700",
		16#10ca# => X"23a4e500",
		16#10cb# => X"6ff0dff8",
		16#10cc# => X"93d59700",
		16#10cd# => X"13074000",
		16#10ce# => X"6368b704",
		16#10cf# => X"13d76700",
		16#10d0# => X"13078703",
		16#10d1# => X"93051700",
		16#10d2# => X"93953500",
		16#10d3# => X"b305b600",
		16#10d4# => X"138585ff",
		16#10d5# => X"83a50500",
		16#10d6# => X"6314b508",
		16#10d7# => X"93071000",
		16#10d8# => X"13572740",
		16#10d9# => X"3397e700",
		16#10da# => X"83274600",
		16#10db# => X"3367f700",
		16#10dc# => X"2322e600",
		16#10dd# => X"23a6a600",
		16#10de# => X"23a4b600",
		16#10df# => X"2324d500",
		16#10e0# => X"23a6d500",
		16#10e1# => X"6ff0dfea",
		16#10e2# => X"13074001",
		16#10e3# => X"6366b700",
		16#10e4# => X"1387b505",
		16#10e5# => X"6ff01ffb",
		16#10e6# => X"13074005",
		16#10e7# => X"6368b700",
		16#10e8# => X"13d7c700",
		16#10e9# => X"1307e706",
		16#10ea# => X"6ff0dff9",
		16#10eb# => X"13074015",
		16#10ec# => X"6368b700",
		16#10ed# => X"13d7f700",
		16#10ee# => X"13077707",
		16#10ef# => X"6ff09ff8",
		16#10f0# => X"13054055",
		16#10f1# => X"1307e007",
		16#10f2# => X"e36eb5f6",
		16#10f3# => X"13d72701",
		16#10f4# => X"1307c707",
		16#10f5# => X"6ff01ff7",
		16#10f6# => X"83a58500",
		16#10f7# => X"6308b500",
		16#10f8# => X"03a74500",
		16#10f9# => X"1377c7ff",
		16#10fa# => X"e3e8e7fe",
		16#10fb# => X"03a5c500",
		16#10fc# => X"6ff05ff8",
		16#10fd# => X"67800000",
		16#10fe# => X"83278600",
		16#10ff# => X"63980700",
		16#1100# => X"93070000",
		16#1101# => X"13850700",
		16#1102# => X"67800000",
		16#1103# => X"83d7c500",
		16#1104# => X"130101fc",
		16#1105# => X"232c8102",
		16#1106# => X"23282103",
		16#1107# => X"23206103",
		16#1108# => X"232e1102",
		16#1109# => X"232a9102",
		16#110a# => X"23263103",
		16#110b# => X"23244103",
		16#110c# => X"23225103",
		16#110d# => X"232e7101",
		16#110e# => X"232c8101",
		16#110f# => X"232a9101",
		16#1110# => X"2328a101",
		16#1111# => X"2326b101",
		16#1112# => X"93f78700",
		16#1113# => X"130b0600",
		16#1114# => X"13840500",
		16#1115# => X"13090500",
		16#1116# => X"6382070e",
		16#1117# => X"83a70501",
		16#1118# => X"638e070c",
		16#1119# => X"8357c400",
		16#111a# => X"032a0b00",
		16#111b# => X"13f72700",
		16#111c# => X"631a0716",
		16#111d# => X"93f71700",
		16#111e# => X"930b0000",
		16#111f# => X"638a0720",
		16#1120# => X"13050000",
		16#1121# => X"930a0000",
		16#1122# => X"93090000",
		16#1123# => X"63860936",
		16#1124# => X"63120502",
		16#1125# => X"13860900",
		16#1126# => X"9305a000",
		16#1127# => X"13850a00",
		16#1128# => X"ef20d06d",
		16#1129# => X"938b1900",
		16#112a# => X"63060500",
		16#112b# => X"13051500",
		16#112c# => X"b30b5541",
		16#112d# => X"138c0b00",
		16#112e# => X"63f47901",
		16#112f# => X"138c0900",
		16#1130# => X"03250400",
		16#1131# => X"83270401",
		16#1132# => X"83264401",
		16#1133# => X"63f0a734",
		16#1134# => X"83248400",
		16#1135# => X"b3849600",
		16#1136# => X"63da8433",
		16#1137# => X"93850a00",
		16#1138# => X"13860400",
		16#1139# => X"ef20507a",
		16#113a# => X"83270400",
		16#113b# => X"93050400",
		16#113c# => X"13050900",
		16#113d# => X"b3879700",
		16#113e# => X"2320f400",
		16#113f# => X"eff01f85",
		16#1140# => X"631e0516",
		16#1141# => X"b38b9b40",
		16#1142# => X"13051000",
		16#1143# => X"639a0b00",
		16#1144# => X"93050400",
		16#1145# => X"13050900",
		16#1146# => X"eff05f83",
		16#1147# => X"63100516",
		16#1148# => X"83278b00",
		16#1149# => X"b38a9a00",
		16#114a# => X"b3899940",
		16#114b# => X"b3849740",
		16#114c# => X"23249b00",
		16#114d# => X"e39c04f4",
		16#114e# => X"6f008006",
		16#114f# => X"93050400",
		16#1150# => X"13050900",
		16#1151# => X"eff0cfcc",
		16#1152# => X"9307f0ff",
		16#1153# => X"e30c05f0",
		16#1154# => X"6f004005",
		16#1155# => X"83290a00",
		16#1156# => X"83244a00",
		16#1157# => X"130a8a00",
		16#1158# => X"e38a04fe",
		16#1159# => X"93860400",
		16#115a# => X"63f49a00",
		16#115b# => X"93860a00",
		16#115c# => X"83274402",
		16#115d# => X"8325c401",
		16#115e# => X"13860900",
		16#115f# => X"13050900",
		16#1160# => X"e7800700",
		16#1161# => X"635ca00e",
		16#1162# => X"83278b00",
		16#1163# => X"b389a900",
		16#1164# => X"b384a440",
		16#1165# => X"3385a740",
		16#1166# => X"2324ab00",
		16#1167# => X"e31205fc",
		16#1168# => X"93070000",
		16#1169# => X"8320c103",
		16#116a# => X"03248103",
		16#116b# => X"83244103",
		16#116c# => X"03290103",
		16#116d# => X"8329c102",
		16#116e# => X"032a8102",
		16#116f# => X"832a4102",
		16#1170# => X"032b0102",
		16#1171# => X"832bc101",
		16#1172# => X"032c8101",
		16#1173# => X"832c4101",
		16#1174# => X"032d0101",
		16#1175# => X"832dc100",
		16#1176# => X"13850700",
		16#1177# => X"13010104",
		16#1178# => X"67800000",
		16#1179# => X"b70a0080",
		16#117a# => X"93090000",
		16#117b# => X"93040000",
		16#117c# => X"93ca0ac0",
		16#117d# => X"6ff0dff6",
		16#117e# => X"832b0a00",
		16#117f# => X"83244a00",
		16#1180# => X"130a8a00",
		16#1181# => X"e38a04fe",
		16#1182# => X"8359c400",
		16#1183# => X"832d8400",
		16#1184# => X"03250400",
		16#1185# => X"93f70920",
		16#1186# => X"63840714",
		16#1187# => X"63e0b40d",
		16#1188# => X"93f70948",
		16#1189# => X"638c070a",
		16#118a# => X"832d0401",
		16#118b# => X"93053000",
		16#118c# => X"330db541",
		16#118d# => X"03254401",
		16#118e# => X"efd0907f",
		16#118f# => X"935af501",
		16#1190# => X"b38aaa00",
		16#1191# => X"93071d00",
		16#1192# => X"93da1a40",
		16#1193# => X"b3879700",
		16#1194# => X"63f4fa00",
		16#1195# => X"938a0700",
		16#1196# => X"93f90940",
		16#1197# => X"6388090c",
		16#1198# => X"93850a00",
		16#1199# => X"13050900",
		16#119a# => X"ef200065",
		16#119b# => X"93090500",
		16#119c# => X"631a0502",
		16#119d# => X"9307c000",
		16#119e# => X"2320f900",
		16#119f# => X"8357c400",
		16#11a0# => X"93e70704",
		16#11a1# => X"2316f400",
		16#11a2# => X"9307f0ff",
		16#11a3# => X"6ff09ff1",
		16#11a4# => X"370c0080",
		16#11a5# => X"934cecff",
		16#11a6# => X"93040000",
		16#11a7# => X"134cfcff",
		16#11a8# => X"6ff05ff6",
		16#11a9# => X"83250401",
		16#11aa# => X"13060d00",
		16#11ab# => X"ef20504f",
		16#11ac# => X"8357c400",
		16#11ad# => X"93f7f7b7",
		16#11ae# => X"93e70708",
		16#11af# => X"2316f400",
		16#11b0# => X"23283401",
		16#11b1# => X"232a5401",
		16#11b2# => X"b389a901",
		16#11b3# => X"b38aaa41",
		16#11b4# => X"23203401",
		16#11b5# => X"938d0400",
		16#11b6# => X"23245401",
		16#11b7# => X"93890400",
		16#11b8# => X"63f4b401",
		16#11b9# => X"938d0400",
		16#11ba# => X"03250400",
		16#11bb# => X"13860d00",
		16#11bc# => X"93850b00",
		16#11bd# => X"ef205059",
		16#11be# => X"83278400",
		16#11bf# => X"b387b741",
		16#11c0# => X"2324f400",
		16#11c1# => X"83270400",
		16#11c2# => X"b38db701",
		16#11c3# => X"2320b401",
		16#11c4# => X"83278b00",
		16#11c5# => X"b38b3b01",
		16#11c6# => X"b3843441",
		16#11c7# => X"b3893741",
		16#11c8# => X"23243b01",
		16#11c9# => X"e39009ee",
		16#11ca# => X"6ff09fe7",
		16#11cb# => X"13860a00",
		16#11cc# => X"93850d00",
		16#11cd# => X"13050900",
		16#11ce# => X"ef30905f",
		16#11cf# => X"93090500",
		16#11d0# => X"e31005f8",
		16#11d1# => X"83250401",
		16#11d2# => X"13050900",
		16#11d3# => X"eff01fa5",
		16#11d4# => X"8357c400",
		16#11d5# => X"93f7f7f7",
		16#11d6# => X"2316f400",
		16#11d7# => X"6ff09ff1",
		16#11d8# => X"83270401",
		16#11d9# => X"63e6a700",
		16#11da# => X"83294401",
		16#11db# => X"63f63405",
		16#11dc# => X"93890d00",
		16#11dd# => X"63f4b401",
		16#11de# => X"93890400",
		16#11df# => X"13860900",
		16#11e0# => X"93850b00",
		16#11e1# => X"ef205050",
		16#11e2# => X"83278400",
		16#11e3# => X"03270400",
		16#11e4# => X"b3873741",
		16#11e5# => X"33073701",
		16#11e6# => X"2324f400",
		16#11e7# => X"2320e400",
		16#11e8# => X"e39807f6",
		16#11e9# => X"93050400",
		16#11ea# => X"13050900",
		16#11eb# => X"eff00fda",
		16#11ec# => X"e30005f6",
		16#11ed# => X"6ff09fec",
		16#11ee# => X"13050c00",
		16#11ef# => X"63e49c00",
		16#11f0# => X"13850400",
		16#11f1# => X"93850900",
		16#11f2# => X"efd0d068",
		16#11f3# => X"93850900",
		16#11f4# => X"efd01066",
		16#11f5# => X"83274402",
		16#11f6# => X"8325c401",
		16#11f7# => X"93060500",
		16#11f8# => X"13860b00",
		16#11f9# => X"13050900",
		16#11fa# => X"e7800700",
		16#11fb# => X"93090500",
		16#11fc# => X"e340a0f2",
		16#11fd# => X"6ff09fe8",
		16#11fe# => X"832a0a00",
		16#11ff# => X"83294a00",
		16#1200# => X"13050000",
		16#1201# => X"130a8a00",
		16#1202# => X"6ff05fc8",
		16#1203# => X"6342dc02",
		16#1204# => X"83274402",
		16#1205# => X"8325c401",
		16#1206# => X"13860a00",
		16#1207# => X"13050900",
		16#1208# => X"e7800700",
		16#1209# => X"93040500",
		16#120a# => X"e34ea0cc",
		16#120b# => X"6ff01fe5",
		16#120c# => X"13060c00",
		16#120d# => X"93850a00",
		16#120e# => X"ef201045",
		16#120f# => X"83278400",
		16#1210# => X"93040c00",
		16#1211# => X"b3878741",
		16#1212# => X"2324f400",
		16#1213# => X"83270400",
		16#1214# => X"b3878701",
		16#1215# => X"2320f400",
		16#1216# => X"6ff0dfca",
		16#1217# => X"130101fd",
		16#1218# => X"23248102",
		16#1219# => X"23202103",
		16#121a# => X"232c4101",
		16#121b# => X"232a5101",
		16#121c# => X"23261102",
		16#121d# => X"23229102",
		16#121e# => X"232e3101",
		16#121f# => X"1304052e",
		16#1220# => X"13090000",
		16#1221# => X"130a1000",
		16#1222# => X"930af0ff",
		16#1223# => X"63160402",
		16#1224# => X"8320c102",
		16#1225# => X"03248102",
		16#1226# => X"13050900",
		16#1227# => X"83244102",
		16#1228# => X"03290102",
		16#1229# => X"8329c101",
		16#122a# => X"032a8101",
		16#122b# => X"832a4101",
		16#122c# => X"13010103",
		16#122d# => X"67800000",
		16#122e# => X"83248400",
		16#122f# => X"83294400",
		16#1230# => X"9389f9ff",
		16#1231# => X"63d60900",
		16#1232# => X"03240400",
		16#1233# => X"6ff01ffc",
		16#1234# => X"83d7c400",
		16#1235# => X"6370fa02",
		16#1236# => X"8397e400",
		16#1237# => X"638c5701",
		16#1238# => X"13850400",
		16#1239# => X"2326b100",
		16#123a# => X"e7800500",
		16#123b# => X"8325c100",
		16#123c# => X"3369a900",
		16#123d# => X"93848406",
		16#123e# => X"6ff09ffc",
		16#123f# => X"130101fd",
		16#1240# => X"23248102",
		16#1241# => X"23202103",
		16#1242# => X"232c4101",
		16#1243# => X"232a5101",
		16#1244# => X"23286101",
		16#1245# => X"23267101",
		16#1246# => X"23261102",
		16#1247# => X"23229102",
		16#1248# => X"232e3101",
		16#1249# => X"130a0500",
		16#124a# => X"938a0500",
		16#124b# => X"1304052e",
		16#124c# => X"13090000",
		16#124d# => X"130b1000",
		16#124e# => X"930bf0ff",
		16#124f# => X"631a0402",
		16#1250# => X"8320c102",
		16#1251# => X"03248102",
		16#1252# => X"13050900",
		16#1253# => X"83244102",
		16#1254# => X"03290102",
		16#1255# => X"8329c101",
		16#1256# => X"032a8101",
		16#1257# => X"832a4101",
		16#1258# => X"032b0101",
		16#1259# => X"832bc100",
		16#125a# => X"13010103",
		16#125b# => X"67800000",
		16#125c# => X"83248400",
		16#125d# => X"83294400",
		16#125e# => X"9389f9ff",
		16#125f# => X"63d60900",
		16#1260# => X"03240400",
		16#1261# => X"6ff09ffb",
		16#1262# => X"83d7c400",
		16#1263# => X"637efb00",
		16#1264# => X"8397e400",
		16#1265# => X"638a7701",
		16#1266# => X"93850400",
		16#1267# => X"13050a00",
		16#1268# => X"e7800a00",
		16#1269# => X"3369a900",
		16#126a# => X"93848406",
		16#126b# => X"6ff0dffc",
		16#126c# => X"93074501",
		16#126d# => X"13052500",
		16#126e# => X"231f05fe",
		16#126f# => X"e31cf5fe",
		16#1270# => X"67800000",
		16#1271# => X"93074501",
		16#1272# => X"13052500",
		16#1273# => X"0357e5ff",
		16#1274# => X"93852500",
		16#1275# => X"239fe5fe",
		16#1276# => X"e398a7fe",
		16#1277# => X"67800000",
		16#1278# => X"9307a501",
		16#1279# => X"13052500",
		16#127a# => X"231f05fe",
		16#127b# => X"e31cf5fe",
		16#127c# => X"67800000",
		16#127d# => X"13078501",
		16#127e# => X"93870500",
		16#127f# => X"13052500",
		16#1280# => X"8356e5ff",
		16#1281# => X"93872700",
		16#1282# => X"239fd7fe",
		16#1283# => X"e318a7fe",
		16#1284# => X"239c0500",
		16#1285# => X"67800000",
		16#1286# => X"93074500",
		16#1287# => X"93854500",
		16#1288# => X"1305a501",
		16#1289# => X"93872700",
		16#128a# => X"93852500",
		16#128b# => X"83d6e7ff",
		16#128c# => X"03d7e5ff",
		16#128d# => X"6398e600",
		16#128e# => X"e316f5fe",
		16#128f# => X"13050000",
		16#1290# => X"67800000",
		16#1291# => X"13051000",
		16#1292# => X"6364d700",
		16#1293# => X"1305f0ff",
		16#1294# => X"67800000",
		16#1295# => X"93064500",
		16#1296# => X"93070000",
		16#1297# => X"1305a501",
		16#1298# => X"3786ffff",
		16#1299# => X"03d70600",
		16#129a# => X"93751700",
		16#129b# => X"63840500",
		16#129c# => X"93e71700",
		16#129d# => X"93f52700",
		16#129e# => X"13571700",
		16#129f# => X"63900502",
		16#12a0# => X"93971700",
		16#12a1# => X"2390e600",
		16#12a2# => X"93970701",
		16#12a3# => X"93862600",
		16#12a4# => X"93d70701",
		16#12a5# => X"e318d5fc",
		16#12a6# => X"67800000",
		16#12a7# => X"3367c700",
		16#12a8# => X"6ff01ffe",
		16#12a9# => X"93066501",
		16#12aa# => X"13070000",
		16#12ab# => X"83d72600",
		16#12ac# => X"13960701",
		16#12ad# => X"13560641",
		16#12ae# => X"63540600",
		16#12af# => X"13671700",
		16#12b0# => X"93971700",
		16#12b1# => X"93970701",
		16#12b2# => X"13762700",
		16#12b3# => X"93d70701",
		16#12b4# => X"63100602",
		16#12b5# => X"13171700",
		16#12b6# => X"2391f600",
		16#12b7# => X"13170701",
		16#12b8# => X"9386e6ff",
		16#12b9# => X"13570701",
		16#12ba# => X"e312d5fc",
		16#12bb# => X"67800000",
		16#12bc# => X"93e71700",
		16#12bd# => X"6ff01ffe",
		16#12be# => X"93074500",
		16#12bf# => X"13070000",
		16#12c0# => X"1305a501",
		16#12c1# => X"83d60700",
		16#12c2# => X"93872700",
		16#12c3# => X"13d68600",
		16#12c4# => X"3367c700",
		16#12c5# => X"239fe7fe",
		16#12c6# => X"13978600",
		16#12c7# => X"13170701",
		16#12c8# => X"13570701",
		16#12c9# => X"e310f5fe",
		16#12ca# => X"67800000",
		16#12cb# => X"93076501",
		16#12cc# => X"13070000",
		16#12cd# => X"83d62700",
		16#12ce# => X"9387e7ff",
		16#12cf# => X"13968600",
		16#12d0# => X"3367c700",
		16#12d1# => X"2392e700",
		16#12d2# => X"13d78600",
		16#12d3# => X"e314f5fe",
		16#12d4# => X"67800000",
		16#12d5# => X"93074500",
		16#12d6# => X"13078501",
		16#12d7# => X"93872700",
		16#12d8# => X"83d60700",
		16#12d9# => X"239fd7fe",
		16#12da# => X"e31af7fe",
		16#12db# => X"231c0500",
		16#12dc# => X"67800000",
		16#12dd# => X"93078501",
		16#12de# => X"1307a501",
		16#12df# => X"93064500",
		16#12e0# => X"9387e7ff",
		16#12e1# => X"03d60700",
		16#12e2# => X"1307e7ff",
		16#12e3# => X"2310c700",
		16#12e4# => X"e398f6fe",
		16#12e5# => X"23120500",
		16#12e6# => X"67800000",
		16#12e7# => X"93858501",
		16#12e8# => X"13076501",
		16#12e9# => X"93060000",
		16#12ea# => X"83572700",
		16#12eb# => X"03d60500",
		16#12ec# => X"1307e7ff",
		16#12ed# => X"9385e5ff",
		16#12ee# => X"b387c700",
		16#12ef# => X"b387d700",
		16#12f0# => X"2391f500",
		16#12f1# => X"93d70701",
		16#12f2# => X"93f61700",
		16#12f3# => X"e31ee5fc",
		16#12f4# => X"67800000",
		16#12f5# => X"93858501",
		16#12f6# => X"13076501",
		16#12f7# => X"93060000",
		16#12f8# => X"83d70500",
		16#12f9# => X"03562700",
		16#12fa# => X"1307e7ff",
		16#12fb# => X"9385e5ff",
		16#12fc# => X"b387c740",
		16#12fd# => X"b387d740",
		16#12fe# => X"2391f500",
		16#12ff# => X"93d70701",
		16#1300# => X"93f61700",
		16#1301# => X"e31ee5fc",
		16#1302# => X"67800000",
		16#1303# => X"130101fb",
		16#1304# => X"232e3103",
		16#1305# => X"b7090100",
		16#1306# => X"23248104",
		16#1307# => X"23229104",
		16#1308# => X"23202105",
		16#1309# => X"232c4103",
		16#130a# => X"23261104",
		16#130b# => X"130a0500",
		16#130c# => X"23150102",
		16#130d# => X"23160102",
		16#130e# => X"93848501",
		16#130f# => X"13894500",
		16#1310# => X"1304c102",
		16#1311# => X"9389f9ff",
		16#1312# => X"03d50400",
		16#1313# => X"1304e4ff",
		16#1314# => X"9384e4ff",
		16#1315# => X"63180504",
		16#1316# => X"231f04fe",
		16#1317# => X"e31699fe",
		16#1318# => X"93074000",
		16#1319# => X"1307a001",
		16#131a# => X"93054101",
		16#131b# => X"b385f500",
		16#131c# => X"83d50500",
		16#131d# => X"b306f600",
		16#131e# => X"93872700",
		16#131f# => X"2390b600",
		16#1320# => X"e394e7fe",
		16#1321# => X"8320c104",
		16#1322# => X"03248104",
		16#1323# => X"83244104",
		16#1324# => X"03290104",
		16#1325# => X"8329c103",
		16#1326# => X"032a8103",
		16#1327# => X"13010105",
		16#1328# => X"67800000",
		16#1329# => X"93050a00",
		16#132a# => X"2326c100",
		16#132b# => X"efd05018",
		16#132c# => X"03572400",
		16#132d# => X"b3773501",
		16#132e# => X"13550501",
		16#132f# => X"b387e700",
		16#1330# => X"03570400",
		16#1331# => X"2311f400",
		16#1332# => X"93d70701",
		16#1333# => X"3305e500",
		16#1334# => X"3305f500",
		16#1335# => X"2310a400",
		16#1336# => X"13550501",
		16#1337# => X"231fa4fe",
		16#1338# => X"0326c100",
		16#1339# => X"6ff09ff7",
		16#133a# => X"83572501",
		16#133b# => X"93c7f7ff",
		16#133c# => X"13971701",
		16#133d# => X"631c0700",
		16#133e# => X"93072501",
		16#133f# => X"13052500",
		16#1340# => X"0357e5ff",
		16#1341# => X"63180700",
		16#1342# => X"e39aa7fe",
		16#1343# => X"13050000",
		16#1344# => X"67800000",
		16#1345# => X"13051000",
		16#1346# => X"67800000",
		16#1347# => X"130101ff",
		16#1348# => X"23248100",
		16#1349# => X"23261100",
		16#134a# => X"13040500",
		16#134b# => X"eff0dffb",
		16#134c# => X"631e0500",
		16#134d# => X"03152401",
		16#134e# => X"1355f501",
		16#134f# => X"8320c100",
		16#1350# => X"03248100",
		16#1351# => X"13010101",
		16#1352# => X"67800000",
		16#1353# => X"13050000",
		16#1354# => X"6ff0dffe",
		16#1355# => X"83172501",
		16#1356# => X"130101ff",
		16#1357# => X"23261100",
		16#1358# => X"23248100",
		16#1359# => X"23229100",
		16#135a# => X"23202101",
		16#135b# => X"63d80706",
		16#135c# => X"9307f0ff",
		16#135d# => X"2390f500",
		16#135e# => X"03572501",
		16#135f# => X"b7870000",
		16#1360# => X"9387f7ff",
		16#1361# => X"33f7e700",
		16#1362# => X"2391e500",
		16#1363# => X"13090501",
		16#1364# => X"6316f706",
		16#1365# => X"13840500",
		16#1366# => X"93040500",
		16#1367# => X"eff0dff4",
		16#1368# => X"63020504",
		16#1369# => X"93076400",
		16#136a# => X"23120400",
		16#136b# => X"1385c4ff",
		16#136c# => X"1309e9ff",
		16#136d# => X"03572900",
		16#136e# => X"93872700",
		16#136f# => X"239fe7fe",
		16#1370# => X"e318a9fe",
		16#1371# => X"8320c100",
		16#1372# => X"03248100",
		16#1373# => X"83244100",
		16#1374# => X"03290100",
		16#1375# => X"13010101",
		16#1376# => X"67800000",
		16#1377# => X"23900500",
		16#1378# => X"6ff09ff9",
		16#1379# => X"93074400",
		16#137a# => X"9305a401",
		16#137b# => X"93872700",
		16#137c# => X"239f07fe",
		16#137d# => X"e39cb7fe",
		16#137e# => X"6ff0dffc",
		16#137f# => X"93876500",
		16#1380# => X"23920500",
		16#1381# => X"1305e5ff",
		16#1382# => X"1309e9ff",
		16#1383# => X"03572900",
		16#1384# => X"93872700",
		16#1385# => X"239fe7fe",
		16#1386# => X"e318a9fe",
		16#1387# => X"239c0500",
		16#1388# => X"6ff05ffa",
		16#1389# => X"130101fb",
		16#138a# => X"23229104",
		16#138b# => X"23202105",
		16#138c# => X"23261104",
		16#138d# => X"23248104",
		16#138e# => X"13090500",
		16#138f# => X"93840500",
		16#1390# => X"eff09fea",
		16#1391# => X"6310050e",
		16#1392# => X"13850400",
		16#1393# => X"eff0dfe9",
		16#1394# => X"13040500",
		16#1395# => X"6318050c",
		16#1396# => X"93058100",
		16#1397# => X"13050900",
		16#1398# => X"eff05fef",
		16#1399# => X"93054102",
		16#139a# => X"13850400",
		16#139b# => X"eff09fee",
		16#139c# => X"03578100",
		16#139d# => X"83574102",
		16#139e# => X"6380e706",
		16#139f# => X"93072000",
		16#13a0# => X"93068001",
		16#13a1# => X"13068100",
		16#13a2# => X"3306f600",
		16#13a3# => X"03560600",
		16#13a4# => X"631c0602",
		16#13a5# => X"13064102",
		16#13a6# => X"3306f600",
		16#13a7# => X"03560600",
		16#13a8# => X"63140602",
		16#13a9# => X"93872700",
		16#13aa# => X"e39ed7fc",
		16#13ab# => X"13050400",
		16#13ac# => X"8320c104",
		16#13ad# => X"03248104",
		16#13ae# => X"83244104",
		16#13af# => X"03290104",
		16#13b0# => X"13010105",
		16#13b1# => X"67800000",
		16#13b2# => X"13041000",
		16#13b3# => X"e30007fe",
		16#13b4# => X"1304f0ff",
		16#13b5# => X"6ff09ffd",
		16#13b6# => X"13061000",
		16#13b7# => X"63840700",
		16#13b8# => X"1306f0ff",
		16#13b9# => X"93070000",
		16#13ba# => X"93058001",
		16#13bb# => X"13078100",
		16#13bc# => X"3307f700",
		16#13bd# => X"83560700",
		16#13be# => X"13074102",
		16#13bf# => X"3307f700",
		16#13c0# => X"03570700",
		16#13c1# => X"6398e600",
		16#13c2# => X"93872700",
		16#13c3# => X"e390b7fe",
		16#13c4# => X"6ff0dff9",
		16#13c5# => X"13040600",
		16#13c6# => X"e36ad7f8",
		16#13c7# => X"3304c040",
		16#13c8# => X"6ff0dff8",
		16#13c9# => X"1304e0ff",
		16#13ca# => X"6ff05ff8",
		16#13cb# => X"83572501",
		16#13cc# => X"93c7f7ff",
		16#13cd# => X"13971701",
		16#13ce# => X"63100702",
		16#13cf# => X"130101ff",
		16#13d0# => X"23261100",
		16#13d1# => X"eff05fda",
		16#13d2# => X"8320c100",
		16#13d3# => X"13351500",
		16#13d4# => X"13010101",
		16#13d5# => X"67800000",
		16#13d6# => X"13050000",
		16#13d7# => X"67800000",
		16#13d8# => X"93072501",
		16#13d9# => X"13052500",
		16#13da# => X"231f05fe",
		16#13db# => X"e31cf5fe",
		16#13dc# => X"83570500",
		16#13dd# => X"37870000",
		16#13de# => X"1307f7ff",
		16#13df# => X"b3e7e700",
		16#13e0# => X"2310f500",
		16#13e1# => X"67800000",
		16#13e2# => X"130101fe",
		16#13e3# => X"232c8100",
		16#13e4# => X"23282101",
		16#13e5# => X"232e1100",
		16#13e6# => X"232a9100",
		16#13e7# => X"23263101",
		16#13e8# => X"23244101",
		16#13e9# => X"23225101",
		16#13ea# => X"13090500",
		16#13eb# => X"13840500",
		16#13ec# => X"63d20510",
		16#13ed# => X"330ab040",
		16#13ee# => X"93090a00",
		16#13ef# => X"93040000",
		16#13f0# => X"930af000",
		16#13f1# => X"63ce3a03",
		16#13f2# => X"13554a00",
		16#13f3# => X"930500ff",
		16#13f4# => X"efd00066",
		16#13f5# => X"33048540",
		16#13f6# => X"93090400",
		16#13f7# => X"130a7000",
		16#13f8# => X"634c3a03",
		16#13f9# => X"13553400",
		16#13fa# => X"930580ff",
		16#13fb# => X"efd04064",
		16#13fc# => X"33048500",
		16#13fd# => X"631e0402",
		16#13fe# => X"33359000",
		16#13ff# => X"6f004009",
		16#1400# => X"83578901",
		16#1401# => X"13050900",
		16#1402# => X"938909ff",
		16#1403# => X"b3e4f400",
		16#1404# => X"eff05fb6",
		16#1405# => X"6ff01ffb",
		16#1406# => X"83478901",
		16#1407# => X"13050900",
		16#1408# => X"938989ff",
		16#1409# => X"b3e49700",
		16#140a# => X"eff01fad",
		16#140b# => X"6ff05ffb",
		16#140c# => X"83578901",
		16#140d# => X"13050900",
		16#140e# => X"1304f4ff",
		16#140f# => X"93f71700",
		16#1410# => X"b3e49700",
		16#1411# => X"eff01fa1",
		16#1412# => X"6ff0dffa",
		16#1413# => X"13050900",
		16#1414# => X"eff05fb0",
		16#1415# => X"938404ff",
		16#1416# => X"e3ca99fe",
		16#1417# => X"13554400",
		16#1418# => X"930500ff",
		16#1419# => X"efd0c05c",
		16#141a# => X"3304a400",
		16#141b# => X"93040400",
		16#141c# => X"93097000",
		16#141d# => X"63c69904",
		16#141e# => X"13553400",
		16#141f# => X"930580ff",
		16#1420# => X"efd0005b",
		16#1421# => X"3304a400",
		16#1422# => X"63140404",
		16#1423# => X"13050000",
		16#1424# => X"8320c101",
		16#1425# => X"03248101",
		16#1426# => X"83244101",
		16#1427# => X"03290101",
		16#1428# => X"8329c100",
		16#1429# => X"032a8100",
		16#142a# => X"832a4100",
		16#142b# => X"13010102",
		16#142c# => X"67800000",
		16#142d# => X"93840500",
		16#142e# => X"9309f000",
		16#142f# => X"6ff0dff9",
		16#1430# => X"13050900",
		16#1431# => X"eff09fa6",
		16#1432# => X"938484ff",
		16#1433# => X"6ff09ffa",
		16#1434# => X"13050900",
		16#1435# => X"eff01f9d",
		16#1436# => X"1304f4ff",
		16#1437# => X"6ff0dffa",
		16#1438# => X"83574500",
		16#1439# => X"130101ff",
		16#143a# => X"23229100",
		16#143b# => X"23261100",
		16#143c# => X"23248100",
		16#143d# => X"23202101",
		16#143e# => X"93040500",
		16#143f# => X"63920708",
		16#1440# => X"83176500",
		16#1441# => X"13040000",
		16#1442# => X"1309000a",
		16#1443# => X"63d80702",
		16#1444# => X"13050400",
		16#1445# => X"8320c100",
		16#1446# => X"03248100",
		16#1447# => X"83244100",
		16#1448# => X"03290100",
		16#1449# => X"13010101",
		16#144a# => X"67800000",
		16#144b# => X"13850400",
		16#144c# => X"13040401",
		16#144d# => X"eff01fa2",
		16#144e# => X"e30c24fd",
		16#144f# => X"83d76400",
		16#1450# => X"e38607fe",
		16#1451# => X"83d76400",
		16#1452# => X"93f707f0",
		16#1453# => X"63820702",
		16#1454# => X"1309000a",
		16#1455# => X"83976400",
		16#1456# => X"e3cc07fa",
		16#1457# => X"13850400",
		16#1458# => X"13041400",
		16#1459# => X"eff01f94",
		16#145a# => X"e35689fe",
		16#145b# => X"6ff05ffa",
		16#145c# => X"13850400",
		16#145d# => X"eff09f9b",
		16#145e# => X"13048400",
		16#145f# => X"6ff09ffc",
		16#1460# => X"93f707f0",
		16#1461# => X"13040000",
		16#1462# => X"63860700",
		16#1463# => X"eff0df96",
		16#1464# => X"130480ff",
		16#1465# => X"130900f7",
		16#1466# => X"6f004001",
		16#1467# => X"13850400",
		16#1468# => X"1304f4ff",
		16#1469# => X"eff01f8b",
		16#146a# => X"e34424f7",
		16#146b# => X"83d74400",
		16#146c# => X"e39607fe",
		16#146d# => X"6ff0dff5",
		16#146e# => X"93070501",
		16#146f# => X"13052500",
		16#1470# => X"231f05fe",
		16#1471# => X"e31cf5fe",
		16#1472# => X"b7c7ffff",
		16#1473# => X"2310f500",
		16#1474# => X"b787ffff",
		16#1475# => X"93c7f7ff",
		16#1476# => X"2311f500",
		16#1477# => X"67800000",
		16#1478# => X"13070500",
		16#1479# => X"83560700",
		16#147a# => X"13850500",
		16#147b# => X"83572700",
		16#147c# => X"63860600",
		16#147d# => X"b786ffff",
		16#147e# => X"b3e7d700",
		16#147f# => X"2319f500",
		16#1480# => X"03562700",
		16#1481# => X"b7860000",
		16#1482# => X"9386f6ff",
		16#1483# => X"93076700",
		16#1484# => X"631ed600",
		16#1485# => X"1307a701",
		16#1486# => X"83d60700",
		16#1487# => X"63980602",
		16#1488# => X"93872700",
		16#1489# => X"e39ae7fe",
		16#148a# => X"6ff09fd3",
		16#148b# => X"13050501",
		16#148c# => X"13078701",
		16#148d# => X"93872700",
		16#148e# => X"83d6e7ff",
		16#148f# => X"1305e5ff",
		16#1490# => X"2311d500",
		16#1491# => X"e398e7fe",
		16#1492# => X"67800000",
		16#1493# => X"6ff0dff6",
		16#1494# => X"130101fd",
		16#1495# => X"23229102",
		16#1496# => X"93040500",
		16#1497# => X"13054100",
		16#1498# => X"23248102",
		16#1499# => X"23261102",
		16#149a# => X"13840500",
		16#149b# => X"eff04ff7",
		16#149c# => X"03d7e400",
		16#149d# => X"93170701",
		16#149e# => X"93d70741",
		16#149f# => X"63c20704",
		16#14a0# => X"23120100",
		16#14a1# => X"b7860000",
		16#14a2# => X"9386f6ff",
		16#14a3# => X"3377d700",
		16#14a4# => X"9387e400",
		16#14a5# => X"631cd706",
		16#14a6# => X"13870400",
		16#14a7# => X"83560700",
		16#14a8# => X"63860602",
		16#14a9# => X"13050400",
		16#14aa# => X"eff01ff1",
		16#14ab# => X"8320c102",
		16#14ac# => X"03248102",
		16#14ad# => X"83244102",
		16#14ae# => X"13010103",
		16#14af# => X"67800000",
		16#14b0# => X"9307f0ff",
		16#14b1# => X"2312f100",
		16#14b2# => X"6ff0dffb",
		16#14b3# => X"13072700",
		16#14b4# => X"e396e7fc",
		16#14b5# => X"13050400",
		16#14b6# => X"eff08fed",
		16#14b7# => X"13050400",
		16#14b8# => X"eff01fc8",
		16#14b9# => X"8397e400",
		16#14ba# => X"e3d207fc",
		16#14bb# => X"13050400",
		16#14bc# => X"eff09f9f",
		16#14bd# => X"e31c05fa",
		16#14be# => X"83572401",
		16#14bf# => X"3787ffff",
		16#14c0# => X"b3c7e700",
		16#14c1# => X"2319f400",
		16#14c2# => X"6ff05ffa",
		16#14c3# => X"2313e100",
		16#14c4# => X"93064100",
		16#14c5# => X"9387e7ff",
		16#14c6# => X"03d60700",
		16#14c7# => X"93862600",
		16#14c8# => X"2392c600",
		16#14c9# => X"e398f4fe",
		16#14ca# => X"631c0700",
		16#14cb# => X"23140100",
		16#14cc# => X"93050400",
		16#14cd# => X"13054100",
		16#14ce# => X"eff09fea",
		16#14cf# => X"6ff01ff7",
		16#14d0# => X"93071000",
		16#14d1# => X"9305f0ff",
		16#14d2# => X"13054100",
		16#14d3# => X"2314f100",
		16#14d4# => X"eff09fc3",
		16#14d5# => X"6ff0dffd",
		16#14d6# => X"130101fe",
		16#14d7# => X"232c8100",
		16#14d8# => X"232a9100",
		16#14d9# => X"23282101",
		16#14da# => X"23263101",
		16#14db# => X"23244101",
		16#14dc# => X"23225101",
		16#14dd# => X"13890600",
		16#14de# => X"13840700",
		16#14df# => X"232e1100",
		16#14e0# => X"93040500",
		16#14e1# => X"93890500",
		16#14e2# => X"130a0600",
		16#14e3# => X"930a0700",
		16#14e4# => X"eff01fd5",
		16#14e5# => X"93070009",
		16#14e6# => X"3309a940",
		16#14e7# => X"63d4a704",
		16#14e8# => X"b7870000",
		16#14e9# => X"9387e7ff",
		16#14ea# => X"63c6272d",
		16#14eb# => X"93872400",
		16#14ec# => X"9384a401",
		16#14ed# => X"93872700",
		16#14ee# => X"239f07fe",
		16#14ef# => X"e39c97fe",
		16#14f0# => X"8320c101",
		16#14f1# => X"03248101",
		16#14f2# => X"83244101",
		16#14f3# => X"03290101",
		16#14f4# => X"8329c100",
		16#14f5# => X"032a8100",
		16#14f6# => X"832a4100",
		16#14f7# => X"13010102",
		16#14f8# => X"67800000",
		16#14f9# => X"635e0900",
		16#14fa# => X"930700f7",
		16#14fb# => X"634cf912",
		16#14fc# => X"93050900",
		16#14fd# => X"13850400",
		16#14fe# => X"eff01fb9",
		16#14ff# => X"63100514",
		16#1500# => X"63860a22",
		16#1501# => X"03274400",
		16#1502# => X"83270400",
		16#1503# => X"6306f706",
		16#1504# => X"1305a401",
		16#1505# => X"eff0cfdc",
		16#1506# => X"83274400",
		16#1507# => X"13078003",
		16#1508# => X"638ee716",
		16#1509# => X"6340f712",
		16#150a# => X"13078001",
		16#150b# => X"6386e71a",
		16#150c# => X"13075003",
		16#150d# => X"6382e718",
		16#150e# => X"1307c000",
		16#150f# => X"2324e400",
		16#1510# => X"37070180",
		16#1511# => X"1307f7ff",
		16#1512# => X"232ae400",
		16#1513# => X"13071000",
		16#1514# => X"231ce400",
		16#1515# => X"1307b000",
		16#1516# => X"2326e400",
		16#1517# => X"0327c400",
		16#1518# => X"83568401",
		16#1519# => X"13078700",
		16#151a# => X"13171700",
		16#151b# => X"3307e400",
		16#151c# => X"2315d700",
		16#151d# => X"2320f400",
		16#151e# => X"63422003",
		16#151f# => X"03274400",
		16#1520# => X"93070009",
		16#1521# => X"630cf700",
		16#1522# => X"83d78401",
		16#1523# => X"13850400",
		16#1524# => X"93f71700",
		16#1525# => X"b3e9f900",
		16#1526# => X"eff0cfdb",
		16#1527# => X"83268400",
		16#1528# => X"03564401",
		16#1529# => X"83254400",
		16#152a# => X"13971600",
		16#152b# => X"3387e400",
		16#152c# => X"83570700",
		16#152d# => X"b3f7c700",
		16#152e# => X"1306f008",
		16#152f# => X"634ab600",
		16#1530# => X"93861600",
		16#1531# => X"13060700",
		16#1532# => X"9305c000",
		16#1533# => X"63dad510",
		16#1534# => X"83564401",
		16#1535# => X"03560700",
		16#1536# => X"93c6f6ff",
		16#1537# => X"b3f6c600",
		16#1538# => X"2310d700",
		16#1539# => X"03576401",
		16#153a# => X"b376f700",
		16#153b# => X"638a0610",
		16#153c# => X"6312f702",
		16#153d# => X"63940910",
		16#153e# => X"8327c400",
		16#153f# => X"03578401",
		16#1540# => X"93971700",
		16#1541# => X"b387f400",
		16#1542# => X"83d70700",
		16#1543# => X"b3f7e700",
		16#1544# => X"6388070e",
		16#1545# => X"93850400",
		16#1546# => X"1305a401",
		16#1547# => X"eff00fe8",
		16#1548# => X"6f00000e",
		16#1549# => X"93872400",
		16#154a# => X"9384a401",
		16#154b# => X"93872700",
		16#154c# => X"239f07fe",
		16#154d# => X"e39c97fe",
		16#154e# => X"6ff09fe8",
		16#154f# => X"93091000",
		16#1550# => X"6ff01fec",
		16#1551# => X"13070004",
		16#1552# => X"6388e702",
		16#1553# => X"13071007",
		16#1554# => X"e394e7ee",
		16#1555# => X"37870040",
		16#1556# => X"1307f7ff",
		16#1557# => X"9306a000",
		16#1558# => X"232ae400",
		16#1559# => X"2324d400",
		16#155a# => X"3787ffff",
		16#155b# => X"231ce400",
		16#155c# => X"2326d400",
		16#155d# => X"6ff09fee",
		16#155e# => X"13077000",
		16#155f# => X"2324e400",
		16#1560# => X"37070180",
		16#1561# => X"1307f7ff",
		16#1562# => X"232ae400",
		16#1563# => X"13071000",
		16#1564# => X"231ce400",
		16#1565# => X"13076000",
		16#1566# => X"6ff01fec",
		16#1567# => X"93066000",
		16#1568# => X"37078000",
		16#1569# => X"1307f70f",
		16#156a# => X"232ae400",
		16#156b# => X"2324d400",
		16#156c# => X"13070010",
		16#156d# => X"6ff09ffb",
		16#156e# => X"37070004",
		16#156f# => X"1307f77f",
		16#1570# => X"93066000",
		16#1571# => X"232ae400",
		16#1572# => X"37170000",
		16#1573# => X"2324d400",
		16#1574# => X"13070780",
		16#1575# => X"6ff09ff9",
		16#1576# => X"93064000",
		16#1577# => X"6ff05ffc",
		16#1578# => X"03552600",
		16#1579# => X"63040500",
		16#157a# => X"93e71700",
		16#157b# => X"23110600",
		16#157c# => X"93861600",
		16#157d# => X"13062600",
		16#157e# => X"6ff05fed",
		16#157f# => X"e30c0af0",
		16#1580# => X"634c2001",
		16#1581# => X"03274400",
		16#1582# => X"93070009",
		16#1583# => X"6306f700",
		16#1584# => X"13850400",
		16#1585# => X"eff00fc9",
		16#1586# => X"83d74400",
		16#1587# => X"63880700",
		16#1588# => X"13850400",
		16#1589# => X"eff00fc3",
		16#158a# => X"13091900",
		16#158b# => X"b7870000",
		16#158c# => X"239c0400",
		16#158d# => X"9387e7ff",
		16#158e# => X"63d42703",
		16#158f# => X"b787ffff",
		16#1590# => X"93c7f7ff",
		16#1591# => X"2391f400",
		16#1592# => X"93874400",
		16#1593# => X"93848401",
		16#1594# => X"23900700",
		16#1595# => X"93872700",
		16#1596# => X"e39cf4fe",
		16#1597# => X"6ff05fd6",
		16#1598# => X"63560900",
		16#1599# => X"23910400",
		16#159a# => X"6ff09fd5",
		16#159b# => X"23912401",
		16#159c# => X"6ff01fd5",
		16#159d# => X"e3980ad8",
		16#159e# => X"239c0400",
		16#159f# => X"6ff01ffc",
		16#15a0# => X"130101fe",
		16#15a1# => X"23244101",
		16#15a2# => X"035a2500",
		16#15a3# => X"232c8100",
		16#15a4# => X"13840500",
		16#15a5# => X"232e1100",
		16#15a6# => X"232a9100",
		16#15a7# => X"23282101",
		16#15a8# => X"23225101",
		16#15a9# => X"23206101",
		16#15aa# => X"13090600",
		16#15ab# => X"130b4603",
		16#15ac# => X"23263101",
		16#15ad# => X"930a0500",
		16#15ae# => X"eff09fa2",
		16#15af# => X"83542400",
		16#15b0# => X"330aaa40",
		16#15b1# => X"13050400",
		16#15b2# => X"eff09fa1",
		16#15b3# => X"b384a440",
		16#15b4# => X"13050b00",
		16#15b5# => X"eff0cfb0",
		16#15b6# => X"63d24405",
		16#15b7# => X"13050400",
		16#15b8# => X"03248101",
		16#15b9# => X"8320c101",
		16#15ba# => X"8329c100",
		16#15bb# => X"032a8100",
		16#15bc# => X"832a4100",
		16#15bd# => X"032b0100",
		16#15be# => X"93070900",
		16#15bf# => X"93860400",
		16#15c0# => X"03290101",
		16#15c1# => X"83244101",
		16#15c2# => X"13070000",
		16#15c3# => X"13060000",
		16#15c4# => X"93050000",
		16#15c5# => X"13010102",
		16#15c6# => X"6ff01fc4",
		16#15c7# => X"93050400",
		16#15c8# => X"13850a00",
		16#15c9# => X"eff04faf",
		16#15ca# => X"93090000",
		16#15cb# => X"634aa000",
		16#15cc# => X"93050400",
		16#15cd# => X"13850a00",
		16#15ce# => X"eff0cfc9",
		16#15cf# => X"93091000",
		16#15d0# => X"13050b00",
		16#15d1# => X"eff00fb6",
		16#15d2# => X"8357c904",
		16#15d3# => X"13050400",
		16#15d4# => X"9384f4ff",
		16#15d5# => X"b3e9f900",
		16#15d6# => X"23163905",
		16#15d7# => X"eff08fb4",
		16#15d8# => X"6ff09ff7",
		16#15d9# => X"130101f7",
		16#15da# => X"23248108",
		16#15db# => X"23229108",
		16#15dc# => X"23202109",
		16#15dd# => X"232e3107",
		16#15de# => X"23261108",
		16#15df# => X"232c4107",
		16#15e0# => X"232a5107",
		16#15e1# => X"23286107",
		16#15e2# => X"23267107",
		16#15e3# => X"23248107",
		16#15e4# => X"23229107",
		16#15e5# => X"93040500",
		16#15e6# => X"13840500",
		16#15e7# => X"13090600",
		16#15e8# => X"93890600",
		16#15e9# => X"eff04fd4",
		16#15ea# => X"63020504",
		16#15eb# => X"93050900",
		16#15ec# => X"13850400",
		16#15ed# => X"eff00fa1",
		16#15ee# => X"8320c108",
		16#15ef# => X"03248108",
		16#15f0# => X"83244108",
		16#15f1# => X"03290108",
		16#15f2# => X"8329c107",
		16#15f3# => X"032a8107",
		16#15f4# => X"832a4107",
		16#15f5# => X"032b0107",
		16#15f6# => X"832bc106",
		16#15f7# => X"032c8106",
		16#15f8# => X"832c4106",
		16#15f9# => X"13010109",
		16#15fa# => X"67800000",
		16#15fb# => X"13050400",
		16#15fc# => X"eff08fcf",
		16#15fd# => X"63080500",
		16#15fe# => X"93050900",
		16#15ff# => X"13050400",
		16#1600# => X"6ff05ffb",
		16#1601# => X"13850400",
		16#1602# => X"eff04ff2",
		16#1603# => X"63140506",
		16#1604# => X"13050400",
		16#1605# => X"eff08ff1",
		16#1606# => X"630c0500",
		16#1607# => X"b7450110",
		16#1608# => X"938545ce",
		16#1609# => X"13850400",
		16#160a# => X"eff0cfdf",
		16#160b# => X"630e0504",
		16#160c# => X"13850400",
		16#160d# => X"eff08fef",
		16#160e# => X"63180500",
		16#160f# => X"13050400",
		16#1610# => X"eff0cfee",
		16#1611# => X"630c0504",
		16#1612# => X"13850400",
		16#1613# => X"eff00fcd",
		16#1614# => X"93040500",
		16#1615# => X"13050400",
		16#1616# => X"eff04fcc",
		16#1617# => X"638ca402",
		16#1618# => X"b787ffff",
		16#1619# => X"2319f900",
		16#161a# => X"13050900",
		16#161b# => X"eff04fef",
		16#161c# => X"6ff09ff4",
		16#161d# => X"b7450110",
		16#161e# => X"938545ce",
		16#161f# => X"13050400",
		16#1620# => X"eff04fda",
		16#1621# => X"e31605f8",
		16#1622# => X"13050900",
		16#1623# => X"eff0df92",
		16#1624# => X"6ff09ff2",
		16#1625# => X"23190900",
		16#1626# => X"6ff01ffd",
		16#1627# => X"13850400",
		16#1628# => X"9305c100",
		16#1629# => X"eff00fcb",
		16#162a# => X"13050400",
		16#162b# => X"93058102",
		16#162c# => X"eff04fca",
		16#162d# => X"0354e100",
		16#162e# => X"8354a102",
		16#162f# => X"63140402",
		16#1630# => X"93070000",
		16#1631# => X"13076001",
		16#1632# => X"9306c100",
		16#1633# => X"b386f600",
		16#1634# => X"83d62600",
		16#1635# => X"638a0610",
		16#1636# => X"1305c100",
		16#1637# => X"eff05f80",
		16#1638# => X"3304a040",
		16#1639# => X"8357a102",
		16#163a# => X"138c0400",
		16#163b# => X"63920702",
		16#163c# => X"13076001",
		16#163d# => X"93068102",
		16#163e# => X"b386f600",
		16#163f# => X"83d62600",
		16#1640# => X"638e060e",
		16#1641# => X"13058102",
		16#1642# => X"eff08ffd",
		16#1643# => X"338ca440",
		16#1644# => X"83578102",
		16#1645# => X"938b4903",
		16#1646# => X"93848903",
		16#1647# => X"239af902",
		16#1648# => X"8357a102",
		16#1649# => X"138a0b00",
		16#164a# => X"239bf902",
		16#164b# => X"9387e904",
		16#164c# => X"23900400",
		16#164d# => X"93842400",
		16#164e# => X"e39c97fe",
		16#164f# => X"930a0000",
		16#1650# => X"130b0000",
		16#1651# => X"930cc0fe",
		16#1652# => X"9307c100",
		16#1653# => X"b3875701",
		16#1654# => X"03d58701",
		16#1655# => X"630e0500",
		16#1656# => X"93058102",
		16#1657# => X"13064104",
		16#1658# => X"eff0cfaa",
		16#1659# => X"93850b00",
		16#165a# => X"13054104",
		16#165b# => X"eff00fa3",
		16#165c# => X"83d7c904",
		16#165d# => X"13850b00",
		16#165e# => X"938aeaff",
		16#165f# => X"336bfb00",
		16#1660# => X"eff04f9f",
		16#1661# => X"e3929afd",
		16#1662# => X"93078102",
		16#1663# => X"03570a00",
		16#1664# => X"130a2a00",
		16#1665# => X"93872700",
		16#1666# => X"239fe7fe",
		16#1667# => X"e3189afe",
		16#1668# => X"b7c6ffff",
		16#1669# => X"33048401",
		16#166a# => X"93862600",
		16#166b# => X"93870900",
		16#166c# => X"13070004",
		16#166d# => X"b306d400",
		16#166e# => X"13060000",
		16#166f# => X"93050b00",
		16#1670# => X"13058102",
		16#1671# => X"eff05f99",
		16#1672# => X"0357c100",
		16#1673# => X"83578102",
		16#1674# => X"631cf702",
		16#1675# => X"23140102",
		16#1676# => X"93050900",
		16#1677# => X"13058102",
		16#1678# => X"eff01f80",
		16#1679# => X"6ff05fdd",
		16#167a# => X"93872700",
		16#167b# => X"e39ee7ec",
		16#167c# => X"13050900",
		16#167d# => X"efe0dffb",
		16#167e# => X"6ff01fdc",
		16#167f# => X"93872700",
		16#1680# => X"e39ae7ee",
		16#1681# => X"6ff0dffe",
		16#1682# => X"9307f0ff",
		16#1683# => X"2314f102",
		16#1684# => X"6ff09ffc",
		16#1685# => X"130101f7",
		16#1686# => X"23248108",
		16#1687# => X"23229108",
		16#1688# => X"23202109",
		16#1689# => X"232a5107",
		16#168a# => X"23261108",
		16#168b# => X"232e3107",
		16#168c# => X"232c4107",
		16#168d# => X"23286107",
		16#168e# => X"23267107",
		16#168f# => X"23248107",
		16#1690# => X"23229107",
		16#1691# => X"2320a107",
		16#1692# => X"93040500",
		16#1693# => X"13840500",
		16#1694# => X"13090600",
		16#1695# => X"938a0600",
		16#1696# => X"eff00fa9",
		16#1697# => X"63040504",
		16#1698# => X"93050900",
		16#1699# => X"13850400",
		16#169a# => X"efe0dff5",
		16#169b# => X"8320c108",
		16#169c# => X"03248108",
		16#169d# => X"83244108",
		16#169e# => X"03290108",
		16#169f# => X"8329c107",
		16#16a0# => X"032a8107",
		16#16a1# => X"832a4107",
		16#16a2# => X"032b0107",
		16#16a3# => X"832bc106",
		16#16a4# => X"032c8106",
		16#16a5# => X"832c4106",
		16#16a6# => X"032d0106",
		16#16a7# => X"13010109",
		16#16a8# => X"67800000",
		16#16a9# => X"13050400",
		16#16aa# => X"eff00fa4",
		16#16ab# => X"63080500",
		16#16ac# => X"93050900",
		16#16ad# => X"13050400",
		16#16ae# => X"6ff01ffb",
		16#16af# => X"b7490110",
		16#16b0# => X"938549ce",
		16#16b1# => X"13850400",
		16#16b2# => X"eff0cfb5",
		16#16b3# => X"630e051e",
		16#16b4# => X"13850400",
		16#16b5# => X"eff08fc5",
		16#16b6# => X"93090500",
		16#16b7# => X"13050400",
		16#16b8# => X"eff0cfc4",
		16#16b9# => X"63900920",
		16#16ba# => X"63160520",
		16#16bb# => X"13850400",
		16#16bc# => X"9305c100",
		16#16bd# => X"eff00fa6",
		16#16be# => X"13050400",
		16#16bf# => X"93058102",
		16#16c0# => X"eff04fa5",
		16#16c1# => X"8354a102",
		16#16c2# => X"0354e100",
		16#16c3# => X"63940402",
		16#16c4# => X"93070000",
		16#16c5# => X"13076001",
		16#16c6# => X"93068102",
		16#16c7# => X"b386f600",
		16#16c8# => X"83d62600",
		16#16c9# => X"638e061e",
		16#16ca# => X"13058102",
		16#16cb# => X"eff04fdb",
		16#16cc# => X"b304a040",
		16#16cd# => X"8357e100",
		16#16ce# => X"930b0400",
		16#16cf# => X"63920702",
		16#16d0# => X"13076001",
		16#16d1# => X"9306c100",
		16#16d2# => X"b386f600",
		16#16d3# => X"83d62600",
		16#16d4# => X"638e061c",
		16#16d5# => X"1305c100",
		16#16d6# => X"eff08fd8",
		16#16d7# => X"b30ba440",
		16#16d8# => X"83578102",
		16#16d9# => X"0357a102",
		16#16da# => X"93894a03",
		16#16db# => X"239afa02",
		16#16dc# => X"93878a03",
		16#16dd# => X"239bea02",
		16#16de# => X"138a0700",
		16#16df# => X"1387ea04",
		16#16e0# => X"93872700",
		16#16e1# => X"239f07fe",
		16#16e2# => X"e39ce7fe",
		16#16e3# => X"13058102",
		16#16e4# => X"efe05fec",
		16#16e5# => X"035c2101",
		16#16e6# => X"370b0100",
		16#16e7# => X"9305fbff",
		16#16e8# => X"13050c00",
		16#16e9# => X"efc0d028",
		16#16ea# => X"130d0500",
		16#16eb# => X"938ca901",
		16#16ec# => X"130bfbff",
		16#16ed# => X"0355c102",
		16#16ee# => X"8357e102",
		16#16ef# => X"13040b00",
		16#16f0# => X"13150501",
		16#16f1# => X"3305f500",
		16#16f2# => X"636aad00",
		16#16f3# => X"93050c00",
		16#16f4# => X"efc0d028",
		16#16f5# => X"13140501",
		16#16f6# => X"13540401",
		16#16f7# => X"9305c100",
		16#16f8# => X"13050400",
		16#16f9# => X"13064104",
		16#16fa# => X"eff04f82",
		16#16fb# => X"93058102",
		16#16fc# => X"13054104",
		16#16fd# => X"efe05fe2",
		16#16fe# => X"6356a002",
		16#16ff# => X"93054104",
		16#1700# => X"1305c100",
		16#1701# => X"efe01ffd",
		16#1702# => X"93058102",
		16#1703# => X"13054104",
		16#1704# => X"efe09fe0",
		16#1705# => X"634aa012",
		16#1706# => X"1304f4ff",
		16#1707# => X"13140401",
		16#1708# => X"13540401",
		16#1709# => X"93058102",
		16#170a# => X"13054104",
		16#170b# => X"efe09ffa",
		16#170c# => X"13058102",
		16#170d# => X"23108a00",
		16#170e# => X"130a2a00",
		16#170f# => X"efe09ff1",
		16#1710# => X"e31a9af7",
		16#1711# => X"93070000",
		16#1712# => X"93050000",
		16#1713# => X"13076001",
		16#1714# => X"93068102",
		16#1715# => X"b386f600",
		16#1716# => X"83d64600",
		16#1717# => X"93872700",
		16#1718# => X"b3e5d500",
		16#1719# => X"e396e7fe",
		16#171a# => X"b335b000",
		16#171b# => X"93078102",
		16#171c# => X"03d70900",
		16#171d# => X"93892900",
		16#171e# => X"93872700",
		16#171f# => X"239fe7fe",
		16#1720# => X"e3183aff",
		16#1721# => X"b7460000",
		16#1722# => X"b3847441",
		16#1723# => X"9386f6ff",
		16#1724# => X"93870a00",
		16#1725# => X"13070004",
		16#1726# => X"b386d400",
		16#1727# => X"13060000",
		16#1728# => X"13058102",
		16#1729# => X"eff04feb",
		16#172a# => X"0357c100",
		16#172b# => X"83578102",
		16#172c# => X"631af70a",
		16#172d# => X"23140102",
		16#172e# => X"93050900",
		16#172f# => X"13058102",
		16#1730# => X"eff00fd2",
		16#1731# => X"6ff09fda",
		16#1732# => X"938549ce",
		16#1733# => X"13050400",
		16#1734# => X"eff04f95",
		16#1735# => X"e31e05de",
		16#1736# => X"13050900",
		16#1737# => X"eff0cfcd",
		16#1738# => X"6ff0dfd8",
		16#1739# => X"e31a05fe",
		16#173a# => X"13050900",
		16#173b# => X"efe05fcc",
		16#173c# => X"6ff0dfd7",
		16#173d# => X"13850400",
		16#173e# => X"eff04f82",
		16#173f# => X"93040500",
		16#1740# => X"13050400",
		16#1741# => X"eff08f81",
		16#1742# => X"638ca402",
		16#1743# => X"b787ffff",
		16#1744# => X"2319f900",
		16#1745# => X"13050900",
		16#1746# => X"eff08fa4",
		16#1747# => X"6ff01fd5",
		16#1748# => X"93872700",
		16#1749# => X"e39ae7de",
		16#174a# => X"6ff01ffc",
		16#174b# => X"93872700",
		16#174c# => X"e39ae7e0",
		16#174d# => X"0357c100",
		16#174e# => X"83578102",
		16#174f# => X"e318f7fc",
		16#1750# => X"23190900",
		16#1751# => X"6ff01ffd",
		16#1752# => X"1304e4ff",
		16#1753# => X"13140401",
		16#1754# => X"93054104",
		16#1755# => X"1305c100",
		16#1756# => X"13540401",
		16#1757# => X"efe09fe7",
		16#1758# => X"6ff05fec",
		16#1759# => X"9307f0ff",
		16#175a# => X"2314f102",
		16#175b# => X"6ff0dff4",
		16#175c# => X"03ae0500",
		16#175d# => X"03a34500",
		16#175e# => X"83a88500",
		16#175f# => X"83a5c500",
		16#1760# => X"130101e2",
		16#1761# => X"232c811c",
		16#1762# => X"2326b102",
		16#1763# => X"13840700",
		16#1764# => X"83250504",
		16#1765# => X"9307f0ff",
		16#1766# => X"2328f114",
		16#1767# => X"93070009",
		16#1768# => X"2324411d",
		16#1769# => X"2322511d",
		16#176a# => X"232e711b",
		16#176b# => X"232a911b",
		16#176c# => X"232e111c",
		16#176d# => X"232a911c",
		16#176e# => X"2328211d",
		16#176f# => X"2326311d",
		16#1770# => X"2320611d",
		16#1771# => X"232c811b",
		16#1772# => X"2328a11b",
		16#1773# => X"2326b11b",
		16#1774# => X"23260101",
		16#1775# => X"2320c103",
		16#1776# => X"23226102",
		16#1777# => X"23241103",
		16#1778# => X"232af114",
		16#1779# => X"130a0500",
		16#177a# => X"930b0600",
		16#177b# => X"938a0600",
		16#177c# => X"930c0700",
		16#177d# => X"63800502",
		16#177e# => X"83274504",
		16#177f# => X"13071000",
		16#1780# => X"3317f700",
		16#1781# => X"23a2f500",
		16#1782# => X"23a4e500",
		16#1783# => X"ef10d005",
		16#1784# => X"23200a04",
		16#1785# => X"13050102",
		16#1786# => X"93050105",
		16#1787# => X"eff04fc3",
		16#1788# => X"13050105",
		16#1789# => X"efe09fef",
		16#178a# => X"6300050e",
		16#178b# => X"93071000",
		16#178c# => X"2320f400",
		16#178d# => X"93073000",
		16#178e# => X"638cfb0c",
		16#178f# => X"13094001",
		16#1790# => X"638a0b00",
		16#1791# => X"1389faff",
		16#1792# => X"9307a002",
		16#1793# => X"63d42701",
		16#1794# => X"1309a002",
		16#1795# => X"83274115",
		16#1796# => X"13050105",
		16#1797# => X"2328f100",
		16#1798# => X"efe09fe8",
		16#1799# => X"13040500",
		16#179a# => X"6308050a",
		16#179b# => X"b7450110",
		16#179c# => X"93850593",
		16#179d# => X"13054111",
		16#179e# => X"37240000",
		16#179f# => X"ef20d056",
		16#17a0# => X"1304f470",
		16#17a1# => X"83270101",
		16#17a2# => X"13050105",
		16#17a3# => X"23208116",
		16#17a4# => X"232af114",
		16#17a5# => X"eff08f89",
		16#17a6# => X"93094111",
		16#17a7# => X"63180500",
		16#17a8# => X"13050105",
		16#17a9# => X"efe05fe4",
		16#17aa# => X"e30a0518",
		16#17ab# => X"b7270000",
		16#17ac# => X"9387f770",
		16#17ad# => X"23a0fc00",
		16#17ae# => X"93870900",
		16#17af# => X"13060002",
		16#17b0# => X"9306d002",
		16#17b1# => X"03c70700",
		16#17b2# => X"e308c71c",
		16#17b3# => X"e306d71c",
		16#17b4# => X"13840900",
		16#17b5# => X"93871700",
		16#17b6# => X"03c7f7ff",
		16#17b7# => X"93061400",
		16#17b8# => X"a38fe6fe",
		16#17b9# => X"e31e071a",
		16#17ba# => X"13072000",
		16#17bb# => X"93071000",
		16#17bc# => X"6388eb00",
		16#17bd# => X"83270116",
		16#17be# => X"63d42701",
		16#17bf# => X"93070900",
		16#17c0# => X"93060003",
		16#17c1# => X"6f00d01a",
		16#17c2# => X"23200400",
		16#17c3# => X"6ff09ff2",
		16#17c4# => X"13890a00",
		16#17c5# => X"6ff05ff3",
		16#17c6# => X"93070009",
		16#17c7# => X"9305c106",
		16#17c8# => X"13050105",
		16#17c9# => X"232af114",
		16#17ca# => X"efe0dfa9",
		16#17cb# => X"8357e107",
		16#17cc# => X"23220100",
		16#17cd# => X"13970701",
		16#17ce# => X"13570741",
		16#17cf# => X"63500702",
		16#17d0# => X"37870000",
		16#17d1# => X"1307f7ff",
		16#17d2# => X"b3f7e700",
		16#17d3# => X"231ff106",
		16#17d4# => X"b7070100",
		16#17d5# => X"9387f7ff",
		16#17d6# => X"2322f100",
		16#17d7# => X"374b0110",
		16#17d8# => X"13054bce",
		16#17d9# => X"93058108",
		16#17da# => X"13054501",
		16#17db# => X"efe09fa5",
		16#17dc# => X"0357e107",
		16#17dd# => X"b7440110",
		16#17de# => X"93094bce",
		16#17df# => X"938484cf",
		16#17e0# => X"e3100720",
		16#17e1# => X"1307c106",
		16#17e2# => X"93070000",
		16#17e3# => X"93069000",
		16#17e4# => X"03560700",
		16#17e5# => X"63100610",
		16#17e6# => X"93871700",
		16#17e7# => X"13072700",
		16#17e8# => X"e398d7fe",
		16#17e9# => X"9305010c",
		16#17ea# => X"13058108",
		16#17eb# => X"efe09fda",
		16#17ec# => X"93058108",
		16#17ed# => X"1305010c",
		16#17ee# => X"efe0dfa3",
		16#17ef# => X"9305010c",
		16#17f0# => X"1305c106",
		16#17f1# => X"efe01fd9",
		16#17f2# => X"9305c106",
		16#17f3# => X"1305010c",
		16#17f4# => X"efe05fa2",
		16#17f5# => X"13060115",
		16#17f6# => X"9305c106",
		16#17f7# => X"13058108",
		16#17f8# => X"eff00fea",
		16#17f9# => X"8354c119",
		16#17fa# => X"639a0400",
		16#17fb# => X"93054bce",
		16#17fc# => X"1305c106",
		16#17fd# => X"efe01fe3",
		16#17fe# => X"6318056a",
		16#17ff# => X"83274100",
		16#1800# => X"638a076e",
		16#1801# => X"9307d002",
		16#1802# => X"230af110",
		16#1803# => X"93073000",
		16#1804# => X"93090900",
		16#1805# => X"6398fb00",
		16#1806# => X"b3098900",
		16#1807# => X"9307a002",
		16#1808# => X"e3c03719",
		16#1809# => X"9307a000",
		16#180a# => X"639af46c",
		16#180b# => X"93071003",
		16#180c# => X"a30af110",
		16#180d# => X"9307e002",
		16#180e# => X"230bf110",
		16#180f# => X"130c7111",
		16#1810# => X"635a3001",
		16#1811# => X"93070003",
		16#1812# => X"a30bf110",
		16#1813# => X"9389f9ff",
		16#1814# => X"130c8111",
		16#1815# => X"13041400",
		16#1816# => X"63dc096a",
		16#1817# => X"b7450110",
		16#1818# => X"13060400",
		16#1819# => X"93854595",
		16#181a# => X"13050c00",
		16#181b# => X"ef20d037",
		16#181c# => X"6ff05fe1",
		16#181d# => X"b7450110",
		16#181e# => X"93854594",
		16#181f# => X"6ff09fdf",
		16#1820# => X"8317c107",
		16#1821# => X"63c80700",
		16#1822# => X"b7450110",
		16#1823# => X"93850595",
		16#1824# => X"6ff05fde",
		16#1825# => X"9305c106",
		16#1826# => X"13850400",
		16#1827# => X"efe09fd8",
		16#1828# => X"e30205f0",
		16#1829# => X"635a0546",
		16#182a# => X"9305410a",
		16#182b# => X"1305c106",
		16#182c# => X"efe05f91",
		16#182d# => X"b7470000",
		16#182e# => X"9387e708",
		16#182f# => X"231bf10a",
		16#1830# => X"93070001",
		16#1831# => X"2324f100",
		16#1832# => X"b7870000",
		16#1833# => X"9387f7ff",
		16#1834# => X"232af100",
		16#1835# => X"b7c7ffff",
		16#1836# => X"93872700",
		16#1837# => X"130d0000",
		16#1838# => X"232cf100",
		16#1839# => X"b7470110",
		16#183a# => X"9387c7da",
		16#183b# => X"3385a701",
		16#183c# => X"93060115",
		16#183d# => X"13068108",
		16#183e# => X"9305410a",
		16#183f# => X"eff09f91",
		16#1840# => X"13058108",
		16#1841# => X"9305c103",
		16#1842# => X"efe0df8b",
		16#1843# => X"83274101",
		16#1844# => X"035ce104",
		16#1845# => X"03278101",
		16#1846# => X"b377fc00",
		16#1847# => X"3385e700",
		16#1848# => X"634aa004",
		16#1849# => X"1305010c",
		16#184a# => X"efe09f88",
		16#184b# => X"131c0c01",
		16#184c# => X"135c0c41",
		16#184d# => X"63580c10",
		16#184e# => X"93070000",
		16#184f# => X"1307c103",
		16#1850# => X"3307f700",
		16#1851# => X"83560700",
		16#1852# => X"1307010c",
		16#1853# => X"3307f700",
		16#1854# => X"03570700",
		16#1855# => X"638ae63a",
		16#1856# => X"13850400",
		16#1857# => X"efe0dfb8",
		16#1858# => X"63060508",
		16#1859# => X"9305010c",
		16#185a# => X"13850400",
		16#185b# => X"efe09f85",
		16#185c# => X"6f00400d",
		16#185d# => X"93070009",
		16#185e# => X"b38da740",
		16#185f# => X"9305010c",
		16#1860# => X"1305c103",
		16#1861# => X"efe01f84",
		16#1862# => X"635eb00b",
		16#1863# => X"9306010c",
		16#1864# => X"13870d00",
		16#1865# => X"1306f000",
		16#1866# => X"6342e604",
		16#1867# => X"13d54d00",
		16#1868# => X"9307010c",
		16#1869# => X"13171500",
		16#186a# => X"3387e700",
		16#186b# => X"930500ff",
		16#186c# => X"232ee100",
		16#186d# => X"efc0c047",
		16#186e# => X"0327c101",
		16#186f# => X"3305b501",
		16#1870# => X"13151500",
		16#1871# => X"3385a900",
		16#1872# => X"83560700",
		16#1873# => X"8357c512",
		16#1874# => X"b3f7d700",
		16#1875# => X"2310f700",
		16#1876# => X"6ff05ff5",
		16#1877# => X"23900600",
		16#1878# => X"130707ff",
		16#1879# => X"93862600",
		16#187a# => X"6ff01ffb",
		16#187b# => X"1305010c",
		16#187c# => X"efe09faf",
		16#187d# => X"63080500",
		16#187e# => X"9305010c",
		16#187f# => X"13850500",
		16#1880# => X"6ff0dff6",
		16#1881# => X"13850400",
		16#1882# => X"efe05fd2",
		16#1883# => X"930d0500",
		16#1884# => X"1305010c",
		16#1885# => X"efe09fd1",
		16#1886# => X"130c0500",
		16#1887# => X"638c0d14",
		16#1888# => X"63040512",
		16#1889# => X"13850400",
		16#188a# => X"efe05faf",
		16#188b# => X"130c0500",
		16#188c# => X"1305010c",
		16#188d# => X"efe09fae",
		16#188e# => X"6318ac10",
		16#188f# => X"1305010c",
		16#1890# => X"efe09ff7",
		16#1891# => X"93070000",
		16#1892# => X"13078108",
		16#1893# => X"3307f700",
		16#1894# => X"83560700",
		16#1895# => X"1307010c",
		16#1896# => X"3307f700",
		16#1897# => X"03570700",
		16#1898# => X"6392e602",
		16#1899# => X"93872700",
		16#189a# => X"13072001",
		16#189b# => X"e39ee7fc",
		16#189c# => X"9305410a",
		16#189d# => X"13058108",
		16#189e# => X"efe0cff4",
		16#189f# => X"83278100",
		16#18a0# => X"3304f400",
		16#18a1# => X"83278100",
		16#18a2# => X"130d4d01",
		16#18a3# => X"93d71700",
		16#18a4# => X"2324f100",
		16#18a5# => X"93074006",
		16#18a6# => X"e316fde4",
		16#18a7# => X"8357610b",
		16#18a8# => X"0357e107",
		16#18a9# => X"9305c106",
		16#18aa# => X"1305410a",
		16#18ab# => X"b387e700",
		16#18ac# => X"37c7ffff",
		16#18ad# => X"130727f7",
		16#18ae# => X"b387e700",
		16#18af# => X"231bf10a",
		16#18b0# => X"efe04ff0",
		16#18b1# => X"13850400",
		16#18b2# => X"93058108",
		16#18b3# => X"efe08fef",
		16#18b4# => X"93040000",
		16#18b5# => X"371d0000",
		16#18b6# => X"93898911",
		16#18b7# => X"930d4010",
		16#18b8# => X"b7470110",
		16#18b9# => X"9387c7d0",
		16#18ba# => X"9305410a",
		16#18bb# => X"13850900",
		16#18bc# => X"338c9700",
		16#18bd# => X"efe01fb3",
		16#18be# => X"e346a0ca",
		16#18bf# => X"9305410a",
		16#18c0# => X"13050c00",
		16#18c1# => X"efe01fb2",
		16#18c2# => X"6348a002",
		16#18c3# => X"1306410a",
		16#18c4# => X"93050600",
		16#18c5# => X"93060115",
		16#18c6# => X"13050c00",
		16#18c7# => X"eff08fef",
		16#18c8# => X"13068108",
		16#18c9# => X"93060115",
		16#18ca# => X"93050600",
		16#18cb# => X"13050c00",
		16#18cc# => X"eff04fc3",
		16#18cd# => X"3304a401",
		16#18ce# => X"93844401",
		16#18cf# => X"135d1d00",
		16#18d0# => X"e390b4fb",
		16#18d1# => X"6ff01fc6",
		16#18d2# => X"13850400",
		16#18d3# => X"9305010c",
		16#18d4# => X"efe04fe7",
		16#18d5# => X"1305010c",
		16#18d6# => X"efe01f99",
		16#18d7# => X"e31405ee",
		16#18d8# => X"8357210d",
		16#18d9# => X"3787ffff",
		16#18da# => X"b3c7e700",
		16#18db# => X"2319f10c",
		16#18dc# => X"6ff05fed",
		16#18dd# => X"e31205e8",
		16#18de# => X"9305c10d",
		16#18df# => X"13850400",
		16#18e0# => X"efe05f9d",
		16#18e1# => X"9305810f",
		16#18e2# => X"1305010c",
		16#18e3# => X"efe09f9c",
		16#18e4# => X"0357c10d",
		16#18e5# => X"835da10f",
		16#18e6# => X"8357e10d",
		16#18e7# => X"1347f7ff",
		16#18e8# => X"13170701",
		16#18e9# => X"13570701",
		16#18ea# => X"231ee10c",
		16#18eb# => X"b387b741",
		16#18ec# => X"6358f008",
		16#18ed# => X"93054111",
		16#18ee# => X"1305810f",
		16#18ef# => X"232ef100",
		16#18f0# => X"efe04fe3",
		16#18f1# => X"9305810f",
		16#18f2# => X"1305c10d",
		16#18f3# => X"efe08fe2",
		16#18f4# => X"9305c10d",
		16#18f5# => X"13054111",
		16#18f6# => X"efe0cfe1",
		16#18f7# => X"8327c101",
		16#18f8# => X"835da10f",
		16#18f9# => X"b307f040",
		16#18fa# => X"1307f0f6",
		16#18fb# => X"63cee708",
		16#18fc# => X"93850700",
		16#18fd# => X"1305c10d",
		16#18fe# => X"efe01fb9",
		16#18ff# => X"13080500",
		16#1900# => X"0357c10d",
		16#1901# => X"8357810f",
		16#1902# => X"232e0101",
		16#1903# => X"9305810f",
		16#1904# => X"1305c10d",
		16#1905# => X"6314f70e",
		16#1906# => X"efe04ff8",
		16#1907# => X"0328c101",
		16#1908# => X"93070115",
		16#1909# => X"13070004",
		16#190a# => X"93860d00",
		16#190b# => X"13060c00",
		16#190c# => X"93050800",
		16#190d# => X"1305810f",
		16#190e# => X"efe01ff2",
		16#190f# => X"6f00c004",
		16#1910# => X"e39407fa",
		16#1911# => X"9305810f",
		16#1912# => X"1305c10d",
		16#1913# => X"232ee100",
		16#1914# => X"efe08fdc",
		16#1915# => X"631a0506",
		16#1916# => X"8357810f",
		16#1917# => X"0327c101",
		16#1918# => X"6388e700",
		16#1919# => X"1305010c",
		16#191a# => X"efe08fd4",
		16#191b# => X"6ff09fdd",
		16#191c# => X"63940d02",
		16#191d# => X"0317e10f",
		16#191e# => X"93070000",
		16#191f# => X"63400702",
		16#1920# => X"1305810f",
		16#1921# => X"efe00fe2",
		16#1922# => X"9305010c",
		16#1923# => X"1305810f",
		16#1924# => X"efe01fd5",
		16#1925# => X"6ff01fdb",
		16#1926# => X"93070000",
		16#1927# => X"13076001",
		16#1928# => X"9306810f",
		16#1929# => X"3386f600",
		16#192a# => X"03562600",
		16#192b# => X"63080600",
		16#192c# => X"938d1d00",
		16#192d# => X"231db10f",
		16#192e# => X"6ff01ffd",
		16#192f# => X"93872700",
		16#1930# => X"e390e7fe",
		16#1931# => X"6ff01fff",
		16#1932# => X"13080000",
		16#1933# => X"e35aa0f2",
		16#1934# => X"93054111",
		16#1935# => X"1305810f",
		16#1936# => X"efe0cfd1",
		16#1937# => X"9305810f",
		16#1938# => X"1305c10d",
		16#1939# => X"efe00fd1",
		16#193a# => X"9305c10d",
		16#193b# => X"13054111",
		16#193c# => X"efe04fd0",
		16#193d# => X"13080c00",
		16#193e# => X"6ff09ff0",
		16#193f# => X"efe08fed",
		16#1940# => X"130c1000",
		16#1941# => X"6ff09ff1",
		16#1942# => X"93872700",
		16#1943# => X"13072001",
		16#1944# => X"e396e7c2",
		16#1945# => X"6ff01fd3",
		16#1946# => X"8357e107",
		16#1947# => X"138c8911",
		16#1948# => X"6388070a",
		16#1949# => X"9305010c",
		16#194a# => X"1305c106",
		16#194b# => X"374c0000",
		16#194c# => X"efe05f82",
		16#194d# => X"130cecff",
		16#194e# => X"130d50fd",
		16#194f# => X"8357810d",
		16#1950# => X"93f77700",
		16#1951# => X"63920706",
		16#1952# => X"9305410a",
		16#1953# => X"1305010c",
		16#1954# => X"efe04fca",
		16#1955# => X"1305410a",
		16#1956# => X"efe0cfcf",
		16#1957# => X"1305410a",
		16#1958# => X"efe04fcf",
		16#1959# => X"9305410a",
		16#195a# => X"1305010c",
		16#195b# => X"efe00fe3",
		16#195c# => X"8357610a",
		16#195d# => X"93873700",
		16#195e# => X"2313f10a",
		16#195f# => X"8357810a",
		16#1960# => X"639a0710",
		16#1961# => X"8357c10b",
		16#1962# => X"63900702",
		16#1963# => X"8357610a",
		16#1964# => X"636cfc00",
		16#1965# => X"9305010c",
		16#1966# => X"1305410a",
		16#1967# => X"1304f4ff",
		16#1968# => X"efe04fc5",
		16#1969# => X"e31ca4f9",
		16#196a# => X"9305c106",
		16#196b# => X"1305010c",
		16#196c# => X"efe01fc3",
		16#196d# => X"6f004002",
		16#196e# => X"1306c106",
		16#196f# => X"93060115",
		16#1970# => X"93050600",
		16#1971# => X"13050c00",
		16#1972# => X"eff0cf99",
		16#1973# => X"1304f4ff",
		16#1974# => X"8317c107",
		16#1975# => X"e3d207fe",
		16#1976# => X"9305010c",
		16#1977# => X"1305c106",
		16#1978# => X"efe04fbe",
		16#1979# => X"93058108",
		16#197a# => X"13850400",
		16#197b# => X"efe08fbd",
		16#197c# => X"93870915",
		16#197d# => X"130d0000",
		16#197e# => X"37fcffff",
		16#197f# => X"938d8902",
		16#1980# => X"2324f100",
		16#1981# => X"83278100",
		16#1982# => X"9305010c",
		16#1983# => X"13850400",
		16#1984# => X"3387a701",
		16#1985# => X"232ae100",
		16#1986# => X"efe0df80",
		16#1987# => X"b389ad01",
		16#1988# => X"03274101",
		16#1989# => X"635ca004",
		16#198a# => X"9305010c",
		16#198b# => X"13050700",
		16#198c# => X"efe04fff",
		16#198d# => X"63480502",
		16#198e# => X"1306010c",
		16#198f# => X"93050600",
		16#1990# => X"93060115",
		16#1991# => X"13850900",
		16#1992# => X"eff0cf91",
		16#1993# => X"13068108",
		16#1994# => X"93060115",
		16#1995# => X"93050600",
		16#1996# => X"13850900",
		16#1997# => X"eff08f90",
		16#1998# => X"33048401",
		16#1999# => X"1357fc01",
		16#199a# => X"330c8701",
		16#199b# => X"130d4d01",
		16#199c# => X"93074010",
		16#199d# => X"135c1c40",
		16#199e# => X"e316fdf8",
		16#199f# => X"13068108",
		16#19a0# => X"93060115",
		16#19a1# => X"93850400",
		16#19a2# => X"13050600",
		16#19a3# => X"eff08fb8",
		16#19a4# => X"6ff05f91",
		16#19a5# => X"1305410a",
		16#19a6# => X"efe0cfbb",
		16#19a7# => X"8357610a",
		16#19a8# => X"93871700",
		16#19a9# => X"6ff05fed",
		16#19aa# => X"1305c106",
		16#19ab# => X"efe08fbf",
		16#19ac# => X"9305410a",
		16#19ad# => X"1305c106",
		16#19ae# => X"efe0cfb3",
		16#19af# => X"1305410a",
		16#19b0# => X"efe04fbe",
		16#19b1# => X"1305410a",
		16#19b2# => X"efe0cfbd",
		16#19b3# => X"9305c106",
		16#19b4# => X"1305410a",
		16#19b5# => X"efe08fcc",
		16#19b6# => X"13060115",
		16#19b7# => X"9305c106",
		16#19b8# => X"13058108",
		16#19b9# => X"efe0dff9",
		16#19ba# => X"1304f4ff",
		16#19bb# => X"8354c119",
		16#19bc# => X"6ff09f8f",
		16#19bd# => X"93070002",
		16#19be# => X"6ff01f91",
		16#19bf# => X"93840403",
		16#19c0# => X"9307e002",
		16#19c1# => X"a30a9110",
		16#19c2# => X"230bf110",
		16#19c3# => X"130c7111",
		16#19c4# => X"93040c00",
		16#19c5# => X"b3878441",
		16#19c6# => X"63d6f904",
		16#19c7# => X"8357c119",
		16#19c8# => X"13074000",
		16#19c9# => X"138cf4ff",
		16#19ca# => X"e35af792",
		16#19cb# => X"13075000",
		16#19cc# => X"6384e708",
		16#19cd# => X"93070c00",
		16#19ce# => X"1306e002",
		16#19cf# => X"93058003",
		16#19d0# => X"93060003",
		16#19d1# => X"9387f7ff",
		16#19d2# => X"03c70700",
		16#19d3# => X"1377f707",
		16#19d4# => X"63d6090a",
		16#19d5# => X"13071003",
		16#19d6# => X"2380e700",
		16#19d7# => X"13041400",
		16#19d8# => X"6ff0df8f",
		16#19d9# => X"1305c106",
		16#19da# => X"efe0cfb3",
		16#19db# => X"9305410a",
		16#19dc# => X"1305c106",
		16#19dd# => X"efe00fa8",
		16#19de# => X"1305410a",
		16#19df# => X"efe08fb2",
		16#19e0# => X"1305410a",
		16#19e1# => X"efe00fb2",
		16#19e2# => X"9305c106",
		16#19e3# => X"1305410a",
		16#19e4# => X"efe0cfc0",
		16#19e5# => X"13060115",
		16#19e6# => X"9305c106",
		16#19e7# => X"13058108",
		16#19e8# => X"efe01fee",
		16#19e9# => X"8347c119",
		16#19ea# => X"93841400",
		16#19eb# => X"93870703",
		16#19ec# => X"a38ff4fe",
		16#19ed# => X"6ff01ff6",
		16#19ee# => X"93058108",
		16#19ef# => X"1305c106",
		16#19f0# => X"efe01fa2",
		16#19f1# => X"93054bce",
		16#19f2# => X"13058108",
		16#19f3# => X"efe08fe5",
		16#19f4# => X"e31205f6",
		16#19f5# => X"e3c40988",
		16#19f6# => X"83c7e4ff",
		16#19f7# => X"938727fd",
		16#19f8# => X"93b71700",
		16#19f9# => X"93c7f7ff",
		16#19fa# => X"b307fc00",
		16#19fb# => X"83c70700",
		16#19fc# => X"93f71700",
		16#19fd# => X"e3840786",
		16#19fe# => X"6ff0dff3",
		16#19ff# => X"6314c702",
		16#1a00# => X"03c7f7ff",
		16#1a01# => X"93068003",
		16#1a02# => X"63e8e600",
		16#1a03# => X"13071700",
		16#1a04# => X"a38fe7fe",
		16#1a05# => X"6ff09f84",
		16#1a06# => X"13041400",
		16#1a07# => X"13071003",
		16#1a08# => X"6ff01fff",
		16#1a09# => X"63e8e500",
		16#1a0a# => X"13071700",
		16#1a0b# => X"2380e700",
		16#1a0c# => X"6ff0df82",
		16#1a0d# => X"2380d700",
		16#1a0e# => X"6ff0dff0",
		16#1a0f# => X"13041400",
		16#1a10# => X"23a08c00",
		16#1a11# => X"93870900",
		16#1a12# => X"9306e002",
		16#1a13# => X"03c70700",
		16#1a14# => X"63160700",
		16#1a15# => X"13075004",
		16#1a16# => X"6f00c002",
		16#1a17# => X"630cd700",
		16#1a18# => X"93871700",
		16#1a19# => X"6ff09ffe",
		16#1a1a# => X"03c71700",
		16#1a1b# => X"93871700",
		16#1a1c# => X"a38fe7fe",
		16#1a1d# => X"03c70700",
		16#1a1e# => X"e31807fe",
		16#1a1f# => X"6ff09ffd",
		16#1a20# => X"9387f7ff",
		16#1a21# => X"83c60700",
		16#1a22# => X"6384e600",
		16#1a23# => X"e3eaf9fe",
		16#1a24# => X"23800700",
		16#1a25# => X"6ff04fe2",
		16#1a26# => X"93871700",
		16#1a27# => X"6ff08fe2",
		16#1a28# => X"13840600",
		16#1a29# => X"6ff00fe3",
		16#1a2a# => X"1304f4ff",
		16#1a2b# => X"23000400",
		16#1a2c# => X"0347f4ff",
		16#1a2d# => X"6316d700",
		16#1a2e# => X"33073441",
		16#1a2f# => X"e3c6e7fe",
		16#1a30# => X"93073000",
		16#1a31# => X"13879a00",
		16#1a32# => X"6394fb02",
		16#1a33# => X"83270116",
		16#1a34# => X"3309f900",
		16#1a35# => X"63580900",
		16#1a36# => X"230a0110",
		16#1a37# => X"23a00c00",
		16#1a38# => X"13840900",
		16#1a39# => X"83a70c00",
		16#1a3a# => X"b38afa00",
		16#1a3b# => X"13873a00",
		16#1a3c# => X"23220a04",
		16#1a3d# => X"93074000",
		16#1a3e# => X"93864701",
		16#1a3f# => X"83254a04",
		16#1a40# => X"6378d706",
		16#1a41# => X"13050a00",
		16#1a42# => X"ef00904b",
		16#1a43# => X"2320aa04",
		16#1a44# => X"93850900",
		16#1a45# => X"93040500",
		16#1a46# => X"ef20c047",
		16#1a47# => X"8327c100",
		16#1a48# => X"63880700",
		16#1a49# => X"33043441",
		16#1a4a# => X"33848400",
		16#1a4b# => X"23a08700",
		16#1a4c# => X"8320c11d",
		16#1a4d# => X"0324811d",
		16#1a4e# => X"13850400",
		16#1a4f# => X"0329011d",
		16#1a50# => X"8324411d",
		16#1a51# => X"8329c11c",
		16#1a52# => X"032a811c",
		16#1a53# => X"832a411c",
		16#1a54# => X"032b011c",
		16#1a55# => X"832bc11b",
		16#1a56# => X"032c811b",
		16#1a57# => X"832c411b",
		16#1a58# => X"032d011b",
		16#1a59# => X"832dc11a",
		16#1a5a# => X"1301011e",
		16#1a5b# => X"67800000",
		16#1a5c# => X"93851500",
		16#1a5d# => X"2322ba04",
		16#1a5e# => X"93971700",
		16#1a5f# => X"6ff0dff7",
		16#1a60# => X"b7870000",
		16#1a61# => X"9387f7ff",
		16#1a62# => X"631cf7ee",
		16#1a63# => X"83274100",
		16#1a64# => X"638207ee",
		16#1a65# => X"b7450110",
		16#1a66# => X"93858593",
		16#1a67# => X"6ff08fcd",
		16#1a68# => X"9307a000",
		16#1a69# => X"9309a002",
		16#1a6a# => X"e39af4d4",
		16#1a6b# => X"93071003",
		16#1a6c# => X"a30af110",
		16#1a6d# => X"9307e002",
		16#1a6e# => X"230bf110",
		16#1a6f# => X"9309a002",
		16#1a70# => X"6ff04fe8",
		16#1a71# => X"83270500",
		16#1a72# => X"130101fc",
		16#1a73# => X"93054101",
		16#1a74# => X"2320f100",
		16#1a75# => X"83274500",
		16#1a76# => X"232e1102",
		16#1a77# => X"2322f100",
		16#1a78# => X"83278500",
		16#1a79# => X"2324f100",
		16#1a7a# => X"8327c500",
		16#1a7b# => X"13050100",
		16#1a7c# => X"2326f100",
		16#1a7d# => X"efe0df85",
		16#1a7e# => X"83576102",
		16#1a7f# => X"13050000",
		16#1a80# => X"93c7f7ff",
		16#1a81# => X"13971701",
		16#1a82# => X"631a0700",
		16#1a83# => X"13054101",
		16#1a84# => X"efe08fad",
		16#1a85# => X"13351500",
		16#1a86# => X"13051500",
		16#1a87# => X"8320c103",
		16#1a88# => X"13010104",
		16#1a89# => X"67800000",
		16#1a8a# => X"1305050f",
		16#1a8b# => X"67800000",
		16#1a8c# => X"83a7c181",
		16#1a8d# => X"03a54703",
		16#1a8e# => X"63160500",
		16#1a8f# => X"37550110",
		16#1a90# => X"130505ca",
		16#1a91# => X"1305050f",
		16#1a92# => X"67800000",
		16#1a93# => X"83a7c181",
		16#1a94# => X"03a54703",
		16#1a95# => X"63160500",
		16#1a96# => X"37550110",
		16#1a97# => X"130505ca",
		16#1a98# => X"1305050f",
		16#1a99# => X"67800000",
		16#1a9a# => X"130101ff",
		16#1a9b# => X"23229100",
		16#1a9c# => X"23261100",
		16#1a9d# => X"23248100",
		16#1a9e# => X"b7440110",
		16#1a9f# => X"63020604",
		16#1aa0# => X"b7450110",
		16#1aa1# => X"9385c595",
		16#1aa2# => X"13050600",
		16#1aa3# => X"13040600",
		16#1aa4# => X"efa09fc0",
		16#1aa5# => X"63060502",
		16#1aa6# => X"93858495",
		16#1aa7# => X"13050400",
		16#1aa8# => X"efa09fbf",
		16#1aa9# => X"630e0500",
		16#1aaa# => X"b7450110",
		16#1aab# => X"938545a7",
		16#1aac# => X"13050400",
		16#1aad# => X"efa05fbe",
		16#1aae# => X"93070000",
		16#1aaf# => X"63140500",
		16#1ab0# => X"93878495",
		16#1ab1# => X"8320c100",
		16#1ab2# => X"03248100",
		16#1ab3# => X"83244100",
		16#1ab4# => X"13850700",
		16#1ab5# => X"13010101",
		16#1ab6# => X"67800000",
		16#1ab7# => X"83a7c181",
		16#1ab8# => X"83a74703",
		16#1ab9# => X"63960700",
		16#1aba# => X"b7570110",
		16#1abb# => X"938707ca",
		16#1abc# => X"03c58712",
		16#1abd# => X"67800000",
		16#1abe# => X"0325c50e",
		16#1abf# => X"67800000",
		16#1ac0# => X"83a7c181",
		16#1ac1# => X"83a74703",
		16#1ac2# => X"63960700",
		16#1ac3# => X"b7570110",
		16#1ac4# => X"938707ca",
		16#1ac5# => X"03a5c70e",
		16#1ac6# => X"67800000",
		16#1ac7# => X"13860500",
		16#1ac8# => X"93050500",
		16#1ac9# => X"03a5c181",
		16#1aca# => X"6ff01ff4",
		16#1acb# => X"130101fa",
		16#1acc# => X"232a9104",
		16#1acd# => X"93840500",
		16#1ace# => X"8395e500",
		16#1acf# => X"232c8104",
		16#1ad0# => X"232e1104",
		16#1ad1# => X"13040600",
		16#1ad2# => X"63de0500",
		16#1ad3# => X"83d7c400",
		16#1ad4# => X"23a00600",
		16#1ad5# => X"93f70708",
		16#1ad6# => X"63980704",
		16#1ad7# => X"93070040",
		16#1ad8# => X"6f00c004",
		16#1ad9# => X"13064101",
		16#1ada# => X"2326d100",
		16#1adb# => X"ef504044",
		16#1adc# => X"8326c100",
		16#1add# => X"e34c05fc",
		16#1ade# => X"03278101",
		16#1adf# => X"b7f70000",
		16#1ae0# => X"37150000",
		16#1ae1# => X"b3f7e700",
		16#1ae2# => X"37e7ffff",
		16#1ae3# => X"b387e700",
		16#1ae4# => X"93b71700",
		16#1ae5# => X"23a0f600",
		16#1ae6# => X"93070040",
		16#1ae7# => X"2320f400",
		16#1ae8# => X"13050580",
		16#1ae9# => X"6f000001",
		16#1aea# => X"93070004",
		16#1aeb# => X"2320f400",
		16#1aec# => X"13050000",
		16#1aed# => X"8320c105",
		16#1aee# => X"03248105",
		16#1aef# => X"83244105",
		16#1af0# => X"13010106",
		16#1af1# => X"67800000",
		16#1af2# => X"83d7c500",
		16#1af3# => X"130101fe",
		16#1af4# => X"232c8100",
		16#1af5# => X"232e1100",
		16#1af6# => X"232a9100",
		16#1af7# => X"23282101",
		16#1af8# => X"93f72700",
		16#1af9# => X"13840500",
		16#1afa# => X"63880702",
		16#1afb# => X"93073404",
		16#1afc# => X"2320f400",
		16#1afd# => X"2328f400",
		16#1afe# => X"93071000",
		16#1aff# => X"232af400",
		16#1b00# => X"8320c101",
		16#1b01# => X"03248101",
		16#1b02# => X"83244101",
		16#1b03# => X"03290101",
		16#1b04# => X"13010102",
		16#1b05# => X"67800000",
		16#1b06# => X"9306c100",
		16#1b07# => X"13068100",
		16#1b08# => X"93040500",
		16#1b09# => X"eff09ff0",
		16#1b0a# => X"83258100",
		16#1b0b# => X"13090500",
		16#1b0c# => X"13850400",
		16#1b0d# => X"ef004008",
		16#1b0e# => X"63100502",
		16#1b0f# => X"8317c400",
		16#1b10# => X"13f70720",
		16#1b11# => X"e31e07fa",
		16#1b12# => X"93f7c7ff",
		16#1b13# => X"93e72700",
		16#1b14# => X"2316f400",
		16#1b15# => X"6ff09ff9",
		16#1b16# => X"b7470010",
		16#1b17# => X"9387c7dc",
		16#1b18# => X"23aef402",
		16#1b19# => X"8357c400",
		16#1b1a# => X"2320a400",
		16#1b1b# => X"2328a400",
		16#1b1c# => X"93e70708",
		16#1b1d# => X"2316f400",
		16#1b1e# => X"83278100",
		16#1b1f# => X"232af400",
		16#1b20# => X"8327c100",
		16#1b21# => X"63820702",
		16#1b22# => X"8315e400",
		16#1b23# => X"13850400",
		16#1b24# => X"ef500037",
		16#1b25# => X"630a0500",
		16#1b26# => X"8357c400",
		16#1b27# => X"93f7c7ff",
		16#1b28# => X"93e71700",
		16#1b29# => X"2316f400",
		16#1b2a# => X"8357c400",
		16#1b2b# => X"3369f900",
		16#1b2c# => X"23162401",
		16#1b2d# => X"6ff0dff4",
		16#1b2e# => X"130101fd",
		16#1b2f# => X"23261102",
		16#1b30# => X"23248102",
		16#1b31# => X"23229102",
		16#1b32# => X"23202103",
		16#1b33# => X"232e3101",
		16#1b34# => X"232c4101",
		16#1b35# => X"232a5101",
		16#1b36# => X"23286101",
		16#1b37# => X"23267101",
		16#1b38# => X"23248101",
		16#1b39# => X"9387b500",
		16#1b3a# => X"13076001",
		16#1b3b# => X"6374f704",
		16#1b3c# => X"93f487ff",
		16#1b3d# => X"63d20404",
		16#1b3e# => X"9307c000",
		16#1b3f# => X"2320f500",
		16#1b40# => X"13050000",
		16#1b41# => X"8320c102",
		16#1b42# => X"03248102",
		16#1b43# => X"83244102",
		16#1b44# => X"03290102",
		16#1b45# => X"8329c101",
		16#1b46# => X"032a8101",
		16#1b47# => X"832a4101",
		16#1b48# => X"032b0101",
		16#1b49# => X"832bc100",
		16#1b4a# => X"032c8100",
		16#1b4b# => X"13010103",
		16#1b4c# => X"67800000",
		16#1b4d# => X"93040001",
		16#1b4e# => X"e3e0b4fc",
		16#1b4f# => X"93090500",
		16#1b50# => X"ef009007",
		16#1b51# => X"37590110",
		16#1b52# => X"9307701f",
		16#1b53# => X"1309c9e0",
		16#1b54# => X"63ea9704",
		16#1b55# => X"13878400",
		16#1b56# => X"3307e900",
		16#1b57# => X"03244700",
		16#1b58# => X"930687ff",
		16#1b59# => X"93d73400",
		16#1b5a# => X"6318d400",
		16#1b5b# => X"0324c700",
		16#1b5c# => X"93872700",
		16#1b5d# => X"63008708",
		16#1b5e# => X"83274400",
		16#1b5f# => X"0327c400",
		16#1b60# => X"83268400",
		16#1b61# => X"93f7c7ff",
		16#1b62# => X"b307f400",
		16#1b63# => X"23a6e600",
		16#1b64# => X"2324d700",
		16#1b65# => X"03a74700",
		16#1b66# => X"13671700",
		16#1b67# => X"23a2e700",
		16#1b68# => X"6f00800a",
		16#1b69# => X"13d79400",
		16#1b6a# => X"9307f003",
		16#1b6b# => X"630a0700",
		16#1b6c# => X"93074000",
		16#1b6d# => X"63e2e70a",
		16#1b6e# => X"93d76400",
		16#1b6f# => X"93878703",
		16#1b70# => X"13871700",
		16#1b71# => X"13173700",
		16#1b72# => X"3307e900",
		16#1b73# => X"03244700",
		16#1b74# => X"930587ff",
		16#1b75# => X"1305f000",
		16#1b76# => X"630cb400",
		16#1b77# => X"03274400",
		16#1b78# => X"1377c7ff",
		16#1b79# => X"33069740",
		16#1b7a# => X"6350c50c",
		16#1b7b# => X"9387f7ff",
		16#1b7c# => X"93871700",
		16#1b7d# => X"03240901",
		16#1b7e# => X"b7550110",
		16#1b7f# => X"93068900",
		16#1b80# => X"938545e1",
		16#1b81# => X"6308d412",
		16#1b82# => X"03274400",
		16#1b83# => X"1306f000",
		16#1b84# => X"1377c7ff",
		16#1b85# => X"33059740",
		16#1b86# => X"635aa60a",
		16#1b87# => X"93e71400",
		16#1b88# => X"2322f400",
		16#1b89# => X"33069400",
		16#1b8a# => X"232ac900",
		16#1b8b# => X"2328c900",
		16#1b8c# => X"93671500",
		16#1b8d# => X"2326d600",
		16#1b8e# => X"2324d600",
		16#1b8f# => X"2322f600",
		16#1b90# => X"3307e400",
		16#1b91# => X"2320a700",
		16#1b92# => X"13850900",
		16#1b93# => X"ef000077",
		16#1b94# => X"13058400",
		16#1b95# => X"6ff01feb",
		16#1b96# => X"93074001",
		16#1b97# => X"63e6e700",
		16#1b98# => X"9307b705",
		16#1b99# => X"6ff0dff5",
		16#1b9a# => X"93074005",
		16#1b9b# => X"63e8e700",
		16#1b9c# => X"93d7c400",
		16#1b9d# => X"9387e706",
		16#1b9e# => X"6ff09ff4",
		16#1b9f# => X"93074015",
		16#1ba0# => X"63e8e700",
		16#1ba1# => X"93d7f400",
		16#1ba2# => X"93877707",
		16#1ba3# => X"6ff05ff3",
		16#1ba4# => X"93064055",
		16#1ba5# => X"9307e007",
		16#1ba6# => X"e3e4e6f2",
		16#1ba7# => X"93d72401",
		16#1ba8# => X"9387c707",
		16#1ba9# => X"6ff0dff1",
		16#1baa# => X"8326c400",
		16#1bab# => X"634c0600",
		16#1bac# => X"83278400",
		16#1bad# => X"23a6d700",
		16#1bae# => X"23a4f600",
		16#1baf# => X"b307e400",
		16#1bb0# => X"6ff05fed",
		16#1bb1# => X"13840600",
		16#1bb2# => X"6ff01ff1",
		16#1bb3# => X"232ad900",
		16#1bb4# => X"2328d900",
		16#1bb5# => X"634c0500",
		16#1bb6# => X"3307e400",
		16#1bb7# => X"83274700",
		16#1bb8# => X"93e71700",
		16#1bb9# => X"2322f700",
		16#1bba# => X"6ff01ff6",
		16#1bbb# => X"9306f01f",
		16#1bbc# => X"03284900",
		16#1bbd# => X"63eae616",
		16#1bbe# => X"13573700",
		16#1bbf# => X"13562740",
		16#1bc0# => X"93061000",
		16#1bc1# => X"13071700",
		16#1bc2# => X"b396c600",
		16#1bc3# => X"13173700",
		16#1bc4# => X"3307e900",
		16#1bc5# => X"b3e60601",
		16#1bc6# => X"2322d900",
		16#1bc7# => X"83260700",
		16#1bc8# => X"130687ff",
		16#1bc9# => X"2326c400",
		16#1bca# => X"2324d400",
		16#1bcb# => X"23208700",
		16#1bcc# => X"23a68600",
		16#1bcd# => X"13d72740",
		16#1bce# => X"13031000",
		16#1bcf# => X"3313e300",
		16#1bd0# => X"03274900",
		16#1bd1# => X"636a6706",
		16#1bd2# => X"b3766700",
		16#1bd3# => X"639c0600",
		16#1bd4# => X"93f7c7ff",
		16#1bd5# => X"13131300",
		16#1bd6# => X"b3766700",
		16#1bd7# => X"93874700",
		16#1bd8# => X"e38a06fe",
		16#1bd9# => X"130ef000",
		16#1bda# => X"93963700",
		16#1bdb# => X"b306d900",
		16#1bdc# => X"13880600",
		16#1bdd# => X"13850700",
		16#1bde# => X"0324c800",
		16#1bdf# => X"6316041b",
		16#1be0# => X"13051500",
		16#1be1# => X"13773500",
		16#1be2# => X"13088800",
		16#1be3# => X"e31607fe",
		16#1be4# => X"13f73700",
		16#1be5# => X"63180720",
		16#1be6# => X"03274900",
		16#1be7# => X"9347f3ff",
		16#1be8# => X"b377f700",
		16#1be9# => X"2322f900",
		16#1bea# => X"03274900",
		16#1beb# => X"13131300",
		16#1bec# => X"63646700",
		16#1bed# => X"631c0320",
		16#1bee# => X"832b8900",
		16#1bef# => X"03a44b00",
		16#1bf0# => X"937ac4ff",
		16#1bf1# => X"63e89a00",
		16#1bf2# => X"33879a40",
		16#1bf3# => X"9307f000",
		16#1bf4# => X"63cee730",
		16#1bf5# => X"03a44184",
		16#1bf6# => X"03a70182",
		16#1bf7# => X"9307f0ff",
		16#1bf8# => X"33848400",
		16#1bf9# => X"6318f71e",
		16#1bfa# => X"13040401",
		16#1bfb# => X"93050400",
		16#1bfc# => X"13850900",
		16#1bfd# => X"ef105029",
		16#1bfe# => X"9307f0ff",
		16#1bff# => X"130b0500",
		16#1c00# => X"630cf526",
		16#1c01# => X"b3875b01",
		16#1c02# => X"6374f500",
		16#1c03# => X"63962b27",
		16#1c04# => X"93860185",
		16#1c05# => X"03a70600",
		16#1c06# => X"138c0185",
		16#1c07# => X"3307e400",
		16#1c08# => X"23a0e600",
		16#1c09# => X"6394671d",
		16#1c0a# => X"93964701",
		16#1c0b# => X"6390061c",
		16#1c0c# => X"83278900",
		16#1c0d# => X"33848a00",
		16#1c0e# => X"13641400",
		16#1c0f# => X"23a28700",
		16#1c10# => X"37570110",
		16#1c11# => X"83270c00",
		16#1c12# => X"83268725",
		16#1c13# => X"63f4f600",
		16#1c14# => X"232cf724",
		16#1c15# => X"37570110",
		16#1c16# => X"83264725",
		16#1c17# => X"63fef620",
		16#1c18# => X"232af724",
		16#1c19# => X"6f004021",
		16#1c1a# => X"13569700",
		16#1c1b# => X"93064000",
		16#1c1c# => X"63e6c604",
		16#1c1d# => X"93566700",
		16#1c1e# => X"93868603",
		16#1c1f# => X"13861600",
		16#1c20# => X"13163600",
		16#1c21# => X"3306c900",
		16#1c22# => X"130586ff",
		16#1c23# => X"03260600",
		16#1c24# => X"6312c508",
		16#1c25# => X"93d62640",
		16#1c26# => X"13071000",
		16#1c27# => X"b316d700",
		16#1c28# => X"b3e60601",
		16#1c29# => X"2322d900",
		16#1c2a# => X"2326a400",
		16#1c2b# => X"2324c400",
		16#1c2c# => X"23248500",
		16#1c2d# => X"23268600",
		16#1c2e# => X"6ff0dfe7",
		16#1c2f# => X"93064001",
		16#1c30# => X"63e6c600",
		16#1c31# => X"9306b605",
		16#1c32# => X"6ff05ffb",
		16#1c33# => X"93064005",
		16#1c34# => X"63e8c600",
		16#1c35# => X"9356c700",
		16#1c36# => X"9386e606",
		16#1c37# => X"6ff01ffa",
		16#1c38# => X"93064015",
		16#1c39# => X"63e8c600",
		16#1c3a# => X"9356f700",
		16#1c3b# => X"93867607",
		16#1c3c# => X"6ff0dff8",
		16#1c3d# => X"13054055",
		16#1c3e# => X"9306e007",
		16#1c3f# => X"e360c5f8",
		16#1c40# => X"93562701",
		16#1c41# => X"9386c607",
		16#1c42# => X"6ff05ff7",
		16#1c43# => X"03268600",
		16#1c44# => X"6308c500",
		16#1c45# => X"83264600",
		16#1c46# => X"93f6c6ff",
		16#1c47# => X"e368d7fe",
		16#1c48# => X"0325c600",
		16#1c49# => X"6ff05ff8",
		16#1c4a# => X"03274400",
		16#1c4b# => X"0326c400",
		16#1c4c# => X"1377c7ff",
		16#1c4d# => X"b3089740",
		16#1c4e# => X"63501e05",
		16#1c4f# => X"93e71400",
		16#1c50# => X"2322f400",
		16#1c51# => X"83278400",
		16#1c52# => X"b3069400",
		16#1c53# => X"3307e400",
		16#1c54# => X"23a6c700",
		16#1c55# => X"2324f600",
		16#1c56# => X"232ad900",
		16#1c57# => X"2328d900",
		16#1c58# => X"93e71800",
		16#1c59# => X"23a6b600",
		16#1c5a# => X"23a4b600",
		16#1c5b# => X"23a2f600",
		16#1c5c# => X"23201701",
		16#1c5d# => X"6ff05fcd",
		16#1c5e# => X"63c20802",
		16#1c5f# => X"3307e400",
		16#1c60# => X"83274700",
		16#1c61# => X"93e71700",
		16#1c62# => X"2322f700",
		16#1c63# => X"83278400",
		16#1c64# => X"23a6c700",
		16#1c65# => X"2324f600",
		16#1c66# => X"6ff01fcb",
		16#1c67# => X"13040600",
		16#1c68# => X"6ff0dfdd",
		16#1c69# => X"138786ff",
		16#1c6a# => X"83a60600",
		16#1c6b# => X"9387f7ff",
		16#1c6c# => X"e380e6de",
		16#1c6d# => X"6ff05fdf",
		16#1c6e# => X"93874700",
		16#1c6f# => X"13131300",
		16#1c70# => X"b3766700",
		16#1c71# => X"e38a06fe",
		16#1c72# => X"6ff01fda",
		16#1c73# => X"93070500",
		16#1c74# => X"6ff01fff",
		16#1c75# => X"b7170000",
		16#1c76# => X"9387f700",
		16#1c77# => X"3304f400",
		16#1c78# => X"b7f7ffff",
		16#1c79# => X"3374f400",
		16#1c7a# => X"6ff05fe0",
		16#1c7b# => X"03a60182",
		16#1c7c# => X"9306f0ff",
		16#1c7d# => X"6316d60a",
		16#1c7e# => X"23a06183",
		16#1c7f# => X"93757b00",
		16#1c80# => X"63880500",
		16#1c81# => X"93078000",
		16#1c82# => X"b385b740",
		16#1c83# => X"330bbb00",
		16#1c84# => X"b7170000",
		16#1c85# => X"b385f500",
		16#1c86# => X"33048b00",
		16#1c87# => X"9387f7ff",
		16#1c88# => X"3374f400",
		16#1c89# => X"338a8540",
		16#1c8a# => X"93050a00",
		16#1c8b# => X"13850900",
		16#1c8c# => X"ef109005",
		16#1c8d# => X"9307f0ff",
		16#1c8e# => X"6316f500",
		16#1c8f# => X"13050b00",
		16#1c90# => X"130a0000",
		16#1c91# => X"83270c00",
		16#1c92# => X"33056541",
		16#1c93# => X"23246901",
		16#1c94# => X"b3874701",
		16#1c95# => X"330a4501",
		16#1c96# => X"136a1a00",
		16#1c97# => X"2320fc00",
		16#1c98# => X"23224b01",
		16#1c99# => X"e38e2bdd",
		16#1c9a# => X"1307f000",
		16#1c9b# => X"63625705",
		16#1c9c# => X"93071000",
		16#1c9d# => X"2322fb00",
		16#1c9e# => X"83278900",
		16#1c9f# => X"83a74700",
		16#1ca0# => X"93f7c7ff",
		16#1ca1# => X"33879740",
		16#1ca2# => X"63e69700",
		16#1ca3# => X"9307f000",
		16#1ca4# => X"63cee704",
		16#1ca5# => X"13850900",
		16#1ca6# => X"ef004032",
		16#1ca7# => X"6ff05fa6",
		16#1ca8# => X"b307fb40",
		16#1ca9# => X"b387e700",
		16#1caa# => X"2320fc00",
		16#1cab# => X"6ff01ff5",
		16#1cac# => X"83a74b00",
		16#1cad# => X"13844aff",
		16#1cae# => X"137484ff",
		16#1caf# => X"93f71700",
		16#1cb0# => X"b3e78700",
		16#1cb1# => X"23a2fb00",
		16#1cb2# => X"93065000",
		16#1cb3# => X"b3878b00",
		16#1cb4# => X"23a2d700",
		16#1cb5# => X"23a4d700",
		16#1cb6# => X"e37487d6",
		16#1cb7# => X"93858b00",
		16#1cb8# => X"13850900",
		16#1cb9# => X"efc09feb",
		16#1cba# => X"6ff09fd5",
		16#1cbb# => X"03248900",
		16#1cbc# => X"93e71400",
		16#1cbd# => X"2322f400",
		16#1cbe# => X"b3079400",
		16#1cbf# => X"2324f900",
		16#1cc0# => X"6ff09fa9",
		16#1cc1# => X"83a7c181",
		16#1cc2# => X"83a74703",
		16#1cc3# => X"63960700",
		16#1cc4# => X"b7570110",
		16#1cc5# => X"938707ca",
		16#1cc6# => X"03a3470e",
		16#1cc7# => X"67000300",
		16#1cc8# => X"639a0502",
		16#1cc9# => X"130101ff",
		16#1cca# => X"9305c100",
		16#1ccb# => X"13050000",
		16#1ccc# => X"630e0600",
		16#1ccd# => X"1305e0ff",
		16#1cce# => X"638a0600",
		16#1ccf# => X"83470600",
		16#1cd0# => X"23a0f500",
		16#1cd1# => X"03450600",
		16#1cd2# => X"3335a000",
		16#1cd3# => X"13010101",
		16#1cd4# => X"67800000",
		16#1cd5# => X"13050000",
		16#1cd6# => X"63000602",
		16#1cd7# => X"1305e0ff",
		16#1cd8# => X"638c0600",
		16#1cd9# => X"83470600",
		16#1cda# => X"23a0f500",
		16#1cdb# => X"03450600",
		16#1cdc# => X"3335a000",
		16#1cdd# => X"67800000",
		16#1cde# => X"67800000",
		16#1cdf# => X"93f5f50f",
		16#1ce0# => X"3306c500",
		16#1ce1# => X"6316c500",
		16#1ce2# => X"13050000",
		16#1ce3# => X"67800000",
		16#1ce4# => X"83470500",
		16#1ce5# => X"e38cb7fe",
		16#1ce6# => X"13051500",
		16#1ce7# => X"6ff09ffe",
		16#1ce8# => X"b3c7a500",
		16#1ce9# => X"93f73700",
		16#1cea# => X"3307c500",
		16#1ceb# => X"63960700",
		16#1cec# => X"93073000",
		16#1ced# => X"63e4c702",
		16#1cee# => X"93070500",
		16#1cef# => X"636ce500",
		16#1cf0# => X"67800000",
		16#1cf1# => X"83c60500",
		16#1cf2# => X"93871700",
		16#1cf3# => X"93851500",
		16#1cf4# => X"a38fd7fe",
		16#1cf5# => X"e3e8e7fe",
		16#1cf6# => X"67800000",
		16#1cf7# => X"93773500",
		16#1cf8# => X"63920708",
		16#1cf9# => X"93070500",
		16#1cfa# => X"9376c7ff",
		16#1cfb# => X"138606fe",
		16#1cfc# => X"63f6c708",
		16#1cfd# => X"83a30500",
		16#1cfe# => X"83a24500",
		16#1cff# => X"83af8500",
		16#1d00# => X"03afc500",
		16#1d01# => X"83ae0501",
		16#1d02# => X"03ae4501",
		16#1d03# => X"03a38501",
		16#1d04# => X"83a8c501",
		16#1d05# => X"93854502",
		16#1d06# => X"93874702",
		16#1d07# => X"03a8c5ff",
		16#1d08# => X"23ae77fc",
		16#1d09# => X"23a057fe",
		16#1d0a# => X"23a2f7ff",
		16#1d0b# => X"23a4e7ff",
		16#1d0c# => X"23a6d7ff",
		16#1d0d# => X"23a8c7ff",
		16#1d0e# => X"23aa67fe",
		16#1d0f# => X"23ac17ff",
		16#1d10# => X"23ae07ff",
		16#1d11# => X"6ff0dffa",
		16#1d12# => X"83c60500",
		16#1d13# => X"93871700",
		16#1d14# => X"93851500",
		16#1d15# => X"a38fd7fe",
		16#1d16# => X"93f63700",
		16#1d17# => X"e39606fe",
		16#1d18# => X"6ff09ff8",
		16#1d19# => X"93070500",
		16#1d1a# => X"6ff01fff",
		16#1d1b# => X"03a60500",
		16#1d1c# => X"93874700",
		16#1d1d# => X"93854500",
		16#1d1e# => X"23aec7fe",
		16#1d1f# => X"e3e8d7fe",
		16#1d20# => X"e3eae7f4",
		16#1d21# => X"67800000",
		16#1d22# => X"3307c500",
		16#1d23# => X"63e8a500",
		16#1d24# => X"93070500",
		16#1d25# => X"639ae702",
		16#1d26# => X"67800000",
		16#1d27# => X"b387c500",
		16#1d28# => X"3306f640",
		16#1d29# => X"e376f5fe",
		16#1d2a# => X"b386c700",
		16#1d2b# => X"63940600",
		16#1d2c# => X"67800000",
		16#1d2d# => X"9387f7ff",
		16#1d2e# => X"83c60700",
		16#1d2f# => X"1307f7ff",
		16#1d30# => X"2300d700",
		16#1d31# => X"6ff05ffe",
		16#1d32# => X"93851500",
		16#1d33# => X"83c6f5ff",
		16#1d34# => X"93871700",
		16#1d35# => X"a38fd7fe",
		16#1d36# => X"6ff0dffb",
		16#1d37# => X"1303f000",
		16#1d38# => X"13070500",
		16#1d39# => X"637ec302",
		16#1d3a# => X"9377f700",
		16#1d3b# => X"6390070a",
		16#1d3c# => X"63920508",
		16#1d3d# => X"937606ff",
		16#1d3e# => X"1376f600",
		16#1d3f# => X"b386e600",
		16#1d40# => X"2320b700",
		16#1d41# => X"2322b700",
		16#1d42# => X"2324b700",
		16#1d43# => X"2326b700",
		16#1d44# => X"13070701",
		16#1d45# => X"e366d7fe",
		16#1d46# => X"63140600",
		16#1d47# => X"67800000",
		16#1d48# => X"b306c340",
		16#1d49# => X"93962600",
		16#1d4a# => X"97020000",
		16#1d4b# => X"b3865600",
		16#1d4c# => X"6780c600",
		16#1d4d# => X"2307b700",
		16#1d4e# => X"a306b700",
		16#1d4f# => X"2306b700",
		16#1d50# => X"a305b700",
		16#1d51# => X"2305b700",
		16#1d52# => X"a304b700",
		16#1d53# => X"2304b700",
		16#1d54# => X"a303b700",
		16#1d55# => X"2303b700",
		16#1d56# => X"a302b700",
		16#1d57# => X"2302b700",
		16#1d58# => X"a301b700",
		16#1d59# => X"2301b700",
		16#1d5a# => X"a300b700",
		16#1d5b# => X"2300b700",
		16#1d5c# => X"67800000",
		16#1d5d# => X"93f5f50f",
		16#1d5e# => X"93968500",
		16#1d5f# => X"b3e5d500",
		16#1d60# => X"93960501",
		16#1d61# => X"b3e5d500",
		16#1d62# => X"6ff0dff6",
		16#1d63# => X"93962700",
		16#1d64# => X"97020000",
		16#1d65# => X"b3865600",
		16#1d66# => X"93820000",
		16#1d67# => X"e78006fa",
		16#1d68# => X"93800200",
		16#1d69# => X"938707ff",
		16#1d6a# => X"3307f740",
		16#1d6b# => X"3306f600",
		16#1d6c# => X"e378c3f6",
		16#1d6d# => X"6ff0dff3",
		16#1d6e# => X"67800000",
		16#1d6f# => X"67800000",
		16#1d70# => X"8327c504",
		16#1d71# => X"130101ff",
		16#1d72# => X"23229100",
		16#1d73# => X"23202101",
		16#1d74# => X"23261100",
		16#1d75# => X"23248100",
		16#1d76# => X"93040500",
		16#1d77# => X"13890500",
		16#1d78# => X"63820704",
		16#1d79# => X"03a7c404",
		16#1d7a# => X"93172900",
		16#1d7b# => X"b307f700",
		16#1d7c# => X"03a50700",
		16#1d7d# => X"63100506",
		16#1d7e# => X"13041000",
		16#1d7f# => X"33142401",
		16#1d80# => X"13065400",
		16#1d81# => X"13162600",
		16#1d82# => X"93051000",
		16#1d83# => X"13850400",
		16#1d84# => X"ef408062",
		16#1d85# => X"63020502",
		16#1d86# => X"23222501",
		16#1d87# => X"23248500",
		16#1d88# => X"6f00c003",
		16#1d89# => X"13061002",
		16#1d8a# => X"93054000",
		16#1d8b# => X"ef40c060",
		16#1d8c# => X"23a6a404",
		16#1d8d# => X"e31805fa",
		16#1d8e# => X"13050000",
		16#1d8f# => X"8320c100",
		16#1d90# => X"03248100",
		16#1d91# => X"83244100",
		16#1d92# => X"03290100",
		16#1d93# => X"13010101",
		16#1d94# => X"67800000",
		16#1d95# => X"03270500",
		16#1d96# => X"23a0e700",
		16#1d97# => X"23280500",
		16#1d98# => X"23260500",
		16#1d99# => X"6ff09ffd",
		16#1d9a# => X"63800502",
		16#1d9b# => X"83a74500",
		16#1d9c# => X"13972700",
		16#1d9d# => X"8327c504",
		16#1d9e# => X"b387e700",
		16#1d9f# => X"03a70700",
		16#1da0# => X"23a0e500",
		16#1da1# => X"23a0b700",
		16#1da2# => X"67800000",
		16#1da3# => X"130101fd",
		16#1da4# => X"23229102",
		16#1da5# => X"83a40501",
		16#1da6# => X"232a5101",
		16#1da7# => X"b70a0100",
		16#1da8# => X"23248102",
		16#1da9# => X"23202103",
		16#1daa# => X"232e3101",
		16#1dab# => X"23286101",
		16#1dac# => X"23267101",
		16#1dad# => X"23248101",
		16#1dae# => X"23261102",
		16#1daf# => X"232c4101",
		16#1db0# => X"23229101",
		16#1db1# => X"130b0500",
		16#1db2# => X"13840500",
		16#1db3# => X"930b0600",
		16#1db4# => X"13890600",
		16#1db5# => X"93894501",
		16#1db6# => X"130c0000",
		16#1db7# => X"938afaff",
		16#1db8# => X"83ac0900",
		16#1db9# => X"93850b00",
		16#1dba# => X"93894900",
		16#1dbb# => X"33f55c01",
		16#1dbc# => X"efa01074",
		16#1dbd# => X"330a2501",
		16#1dbe# => X"93850b00",
		16#1dbf# => X"13d50c01",
		16#1dc0# => X"efa01073",
		16#1dc1# => X"93570a01",
		16#1dc2# => X"3305f500",
		16#1dc3# => X"13590501",
		16#1dc4# => X"337a5a01",
		16#1dc5# => X"13150501",
		16#1dc6# => X"33054501",
		16#1dc7# => X"23aea9fe",
		16#1dc8# => X"130c1c00",
		16#1dc9# => X"e34e9cfa",
		16#1dca# => X"63000906",
		16#1dcb# => X"83278400",
		16#1dcc# => X"63c0f404",
		16#1dcd# => X"83254400",
		16#1dce# => X"13050b00",
		16#1dcf# => X"93851500",
		16#1dd0# => X"eff01fe8",
		16#1dd1# => X"03260401",
		16#1dd2# => X"9305c400",
		16#1dd3# => X"93090500",
		16#1dd4# => X"13062600",
		16#1dd5# => X"13162600",
		16#1dd6# => X"1305c500",
		16#1dd7# => X"eff05fc4",
		16#1dd8# => X"93050400",
		16#1dd9# => X"13050b00",
		16#1dda# => X"eff01ff0",
		16#1ddb# => X"13840900",
		16#1ddc# => X"93874400",
		16#1ddd# => X"93972700",
		16#1dde# => X"b307f400",
		16#1ddf# => X"23a22701",
		16#1de0# => X"93841400",
		16#1de1# => X"23289400",
		16#1de2# => X"13050400",
		16#1de3# => X"8320c102",
		16#1de4# => X"03248102",
		16#1de5# => X"83244102",
		16#1de6# => X"03290102",
		16#1de7# => X"8329c101",
		16#1de8# => X"032a8101",
		16#1de9# => X"832a4101",
		16#1dea# => X"032b0101",
		16#1deb# => X"832bc100",
		16#1dec# => X"032c8100",
		16#1ded# => X"832c4100",
		16#1dee# => X"13010103",
		16#1def# => X"67800000",
		16#1df0# => X"130101fe",
		16#1df1# => X"232c8100",
		16#1df2# => X"23244101",
		16#1df3# => X"13840500",
		16#1df4# => X"130a0500",
		16#1df5# => X"93059000",
		16#1df6# => X"13858600",
		16#1df7# => X"232a9100",
		16#1df8# => X"23282101",
		16#1df9# => X"23225101",
		16#1dfa# => X"232e1100",
		16#1dfb# => X"23263101",
		16#1dfc# => X"93040600",
		16#1dfd# => X"938a0600",
		16#1dfe# => X"13090700",
		16#1dff# => X"efa09065",
		16#1e00# => X"93071000",
		16#1e01# => X"93050000",
		16#1e02# => X"63c2a708",
		16#1e03# => X"13050a00",
		16#1e04# => X"eff01fdb",
		16#1e05# => X"93071000",
		16#1e06# => X"2328f500",
		16#1e07# => X"232a2501",
		16#1e08# => X"93079000",
		16#1e09# => X"63da9706",
		16#1e0a# => X"13099400",
		16#1e0b# => X"93090900",
		16#1e0c# => X"33049400",
		16#1e0d# => X"93891900",
		16#1e0e# => X"83c6f9ff",
		16#1e0f# => X"93050500",
		16#1e10# => X"1306a000",
		16#1e11# => X"938606fd",
		16#1e12# => X"13050a00",
		16#1e13# => X"eff01fe4",
		16#1e14# => X"e39289fe",
		16#1e15# => X"33049900",
		16#1e16# => X"130484ff",
		16#1e17# => X"b3848440",
		16#1e18# => X"b3079400",
		16#1e19# => X"63c05705",
		16#1e1a# => X"8320c101",
		16#1e1b# => X"03248101",
		16#1e1c# => X"83244101",
		16#1e1d# => X"03290101",
		16#1e1e# => X"8329c100",
		16#1e1f# => X"032a8100",
		16#1e20# => X"832a4100",
		16#1e21# => X"13010102",
		16#1e22# => X"67800000",
		16#1e23# => X"93971700",
		16#1e24# => X"93851500",
		16#1e25# => X"6ff05ff7",
		16#1e26# => X"1304a400",
		16#1e27# => X"93049000",
		16#1e28# => X"6ff0dffb",
		16#1e29# => X"13041400",
		16#1e2a# => X"8346f4ff",
		16#1e2b# => X"93050500",
		16#1e2c# => X"1306a000",
		16#1e2d# => X"938606fd",
		16#1e2e# => X"13050a00",
		16#1e2f# => X"eff01fdd",
		16#1e30# => X"6ff01ffa",
		16#1e31# => X"3707ffff",
		16#1e32# => X"3377e500",
		16#1e33# => X"93070500",
		16#1e34# => X"13050000",
		16#1e35# => X"63160700",
		16#1e36# => X"93970701",
		16#1e37# => X"13050001",
		16#1e38# => X"370700ff",
		16#1e39# => X"33f7e700",
		16#1e3a# => X"63160700",
		16#1e3b# => X"13058500",
		16#1e3c# => X"93978700",
		16#1e3d# => X"370700f0",
		16#1e3e# => X"33f7e700",
		16#1e3f# => X"63160700",
		16#1e40# => X"13054500",
		16#1e41# => X"93974700",
		16#1e42# => X"370700c0",
		16#1e43# => X"33f7e700",
		16#1e44# => X"63160700",
		16#1e45# => X"13052500",
		16#1e46# => X"93972700",
		16#1e47# => X"63cc0700",
		16#1e48# => X"13971700",
		16#1e49# => X"63560700",
		16#1e4a# => X"13051500",
		16#1e4b# => X"67800000",
		16#1e4c# => X"13050002",
		16#1e4d# => X"67800000",
		16#1e4e# => X"83270500",
		16#1e4f# => X"13f77700",
		16#1e50# => X"630e0702",
		16#1e51# => X"93f61700",
		16#1e52# => X"13070000",
		16#1e53# => X"639c0600",
		16#1e54# => X"13f72700",
		16#1e55# => X"630c0700",
		16#1e56# => X"93d71700",
		16#1e57# => X"2320f500",
		16#1e58# => X"13071000",
		16#1e59# => X"13050700",
		16#1e5a# => X"67800000",
		16#1e5b# => X"93d72700",
		16#1e5c# => X"2320f500",
		16#1e5d# => X"13072000",
		16#1e5e# => X"6ff0dffe",
		16#1e5f# => X"93960701",
		16#1e60# => X"93d60601",
		16#1e61# => X"13070000",
		16#1e62# => X"63960600",
		16#1e63# => X"93d70701",
		16#1e64# => X"13070001",
		16#1e65# => X"93f6f70f",
		16#1e66# => X"63960600",
		16#1e67# => X"13078700",
		16#1e68# => X"93d78700",
		16#1e69# => X"93f6f700",
		16#1e6a# => X"63960600",
		16#1e6b# => X"13074700",
		16#1e6c# => X"93d74700",
		16#1e6d# => X"93f63700",
		16#1e6e# => X"63960600",
		16#1e6f# => X"13072700",
		16#1e70# => X"93d72700",
		16#1e71# => X"93f61700",
		16#1e72# => X"63980600",
		16#1e73# => X"93d71700",
		16#1e74# => X"63880700",
		16#1e75# => X"13071700",
		16#1e76# => X"2320f500",
		16#1e77# => X"6ff09ff8",
		16#1e78# => X"13070002",
		16#1e79# => X"6ff01ff8",
		16#1e7a# => X"130101ff",
		16#1e7b# => X"23248100",
		16#1e7c# => X"13840500",
		16#1e7d# => X"93051000",
		16#1e7e# => X"23261100",
		16#1e7f# => X"eff05fbc",
		16#1e80# => X"232a8500",
		16#1e81# => X"8320c100",
		16#1e82# => X"03248100",
		16#1e83# => X"13071000",
		16#1e84# => X"2328e500",
		16#1e85# => X"13010101",
		16#1e86# => X"67800000",
		16#1e87# => X"03a70501",
		16#1e88# => X"83270601",
		16#1e89# => X"130101fa",
		16#1e8a# => X"232a9104",
		16#1e8b# => X"23244105",
		16#1e8c# => X"232e1104",
		16#1e8d# => X"232c8104",
		16#1e8e# => X"23282105",
		16#1e8f# => X"23263105",
		16#1e90# => X"23225105",
		16#1e91# => X"23206105",
		16#1e92# => X"232e7103",
		16#1e93# => X"232c8103",
		16#1e94# => X"232a9103",
		16#1e95# => X"2328a103",
		16#1e96# => X"2326b103",
		16#1e97# => X"138a0500",
		16#1e98# => X"93040600",
		16#1e99# => X"6356f700",
		16#1e9a# => X"130a0600",
		16#1e9b# => X"93840500",
		16#1e9c# => X"03290a01",
		16#1e9d# => X"83a90401",
		16#1e9e# => X"83278a00",
		16#1e9f# => X"83254a00",
		16#1ea0# => X"330c3901",
		16#1ea1# => X"63d48701",
		16#1ea2# => X"93851500",
		16#1ea3# => X"eff05fb3",
		16#1ea4# => X"930b4501",
		16#1ea5# => X"931c2c00",
		16#1ea6# => X"130d0500",
		16#1ea7# => X"b38c9b01",
		16#1ea8# => X"93870b00",
		16#1ea9# => X"63e49709",
		16#1eaa# => X"130a4a01",
		16#1eab# => X"13192900",
		16#1eac# => X"b3072a01",
		16#1ead# => X"93844401",
		16#1eae# => X"93992900",
		16#1eaf# => X"2326f100",
		16#1eb0# => X"b70a0100",
		16#1eb1# => X"b3873401",
		16#1eb2# => X"2328f100",
		16#1eb3# => X"938afaff",
		16#1eb4# => X"83270101",
		16#1eb5# => X"63e2f406",
		16#1eb6# => X"63588001",
		16#1eb7# => X"938cccff",
		16#1eb8# => X"83a70c00",
		16#1eb9# => X"638a0718",
		16#1eba# => X"8320c105",
		16#1ebb# => X"03248105",
		16#1ebc# => X"23288d01",
		16#1ebd# => X"13050d00",
		16#1ebe# => X"83244105",
		16#1ebf# => X"03290105",
		16#1ec0# => X"8329c104",
		16#1ec1# => X"032a8104",
		16#1ec2# => X"832a4104",
		16#1ec3# => X"032b0104",
		16#1ec4# => X"832bc103",
		16#1ec5# => X"032c8103",
		16#1ec6# => X"832c4103",
		16#1ec7# => X"032d0103",
		16#1ec8# => X"832dc102",
		16#1ec9# => X"13010106",
		16#1eca# => X"67800000",
		16#1ecb# => X"23a00700",
		16#1ecc# => X"93874700",
		16#1ecd# => X"6ff01ff7",
		16#1ece# => X"83ad0400",
		16#1ecf# => X"b3fd5d01",
		16#1ed0# => X"63880d08",
		16#1ed1# => X"13890b00",
		16#1ed2# => X"13070a00",
		16#1ed3# => X"93090000",
		16#1ed4# => X"03260700",
		16#1ed5# => X"93850d00",
		16#1ed6# => X"03240900",
		16#1ed7# => X"33755601",
		16#1ed8# => X"232ae100",
		16#1ed9# => X"232cc100",
		16#1eda# => X"efa0902c",
		16#1edb# => X"03268101",
		16#1edc# => X"03274101",
		16#1edd# => X"337b5401",
		16#1ede# => X"330b6501",
		16#1edf# => X"13074700",
		16#1ee0# => X"13550601",
		16#1ee1# => X"93850d00",
		16#1ee2# => X"330b3b01",
		16#1ee3# => X"232ae100",
		16#1ee4# => X"232ee100",
		16#1ee5# => X"13540401",
		16#1ee6# => X"efa09029",
		16#1ee7# => X"33058500",
		16#1ee8# => X"13540b01",
		16#1ee9# => X"33058500",
		16#1eea# => X"93590501",
		16#1eeb# => X"337b5b01",
		16#1eec# => X"13150501",
		16#1eed# => X"8327c100",
		16#1eee# => X"03274101",
		16#1eef# => X"13064900",
		16#1ef0# => X"33656501",
		16#1ef1# => X"232ea6fe",
		16#1ef2# => X"6360f70a",
		16#1ef3# => X"23223901",
		16#1ef4# => X"03d92400",
		16#1ef5# => X"63040908",
		16#1ef6# => X"03a40b00",
		16#1ef7# => X"938d0b00",
		16#1ef8# => X"93090a00",
		16#1ef9# => X"93060000",
		16#1efa# => X"03a50900",
		16#1efb# => X"93050900",
		16#1efc# => X"232ad100",
		16#1efd# => X"33755501",
		16#1efe# => X"efa09023",
		16#1eff# => X"03db2d00",
		16#1f00# => X"83264101",
		16#1f01# => X"33745401",
		16#1f02# => X"330b6501",
		16#1f03# => X"330bdb00",
		16#1f04# => X"13150b01",
		16#1f05# => X"33648500",
		16#1f06# => X"23a08d00",
		16#1f07# => X"93894900",
		16#1f08# => X"03d5e9ff",
		16#1f09# => X"13864d00",
		16#1f0a# => X"93050900",
		16#1f0b# => X"232ac100",
		16#1f0c# => X"efa01020",
		16#1f0d# => X"03a44d00",
		16#1f0e# => X"8327c100",
		16#1f0f# => X"135b0b01",
		16#1f10# => X"33745401",
		16#1f11# => X"33048500",
		16#1f12# => X"33046401",
		16#1f13# => X"93560401",
		16#1f14# => X"03264101",
		16#1f15# => X"63eef900",
		16#1f16# => X"23a28d00",
		16#1f17# => X"93844400",
		16#1f18# => X"938b4b00",
		16#1f19# => X"6ff0dfe6",
		16#1f1a# => X"13090600",
		16#1f1b# => X"6ff05fee",
		16#1f1c# => X"930d0600",
		16#1f1d# => X"6ff05ff7",
		16#1f1e# => X"130cfcff",
		16#1f1f# => X"6ff0dfe5",
		16#1f20# => X"130101fe",
		16#1f21# => X"232a9100",
		16#1f22# => X"23282101",
		16#1f23# => X"23263101",
		16#1f24# => X"232e1100",
		16#1f25# => X"232c8100",
		16#1f26# => X"23244101",
		16#1f27# => X"93773600",
		16#1f28# => X"13090500",
		16#1f29# => X"93040600",
		16#1f2a# => X"93890500",
		16#1f2b# => X"63840702",
		16#1f2c# => X"9387f7ff",
		16#1f2d# => X"37470110",
		16#1f2e# => X"130787f3",
		16#1f2f# => X"93972700",
		16#1f30# => X"b307f700",
		16#1f31# => X"03a60700",
		16#1f32# => X"93060000",
		16#1f33# => X"eff01f9c",
		16#1f34# => X"93090500",
		16#1f35# => X"93d42440",
		16#1f36# => X"63800408",
		16#1f37# => X"03248904",
		16#1f38# => X"631e0400",
		16#1f39# => X"93051027",
		16#1f3a# => X"13050900",
		16#1f3b# => X"eff0dfcf",
		16#1f3c# => X"2324a904",
		16#1f3d# => X"13040500",
		16#1f3e# => X"23200500",
		16#1f3f# => X"93f71400",
		16#1f40# => X"63840702",
		16#1f41# => X"93850900",
		16#1f42# => X"13060400",
		16#1f43# => X"13050900",
		16#1f44# => X"eff0dfd0",
		16#1f45# => X"130a0500",
		16#1f46# => X"93850900",
		16#1f47# => X"13050900",
		16#1f48# => X"eff09f94",
		16#1f49# => X"93090a00",
		16#1f4a# => X"93d41440",
		16#1f4b# => X"63860402",
		16#1f4c# => X"03250400",
		16#1f4d# => X"631e0500",
		16#1f4e# => X"13060400",
		16#1f4f# => X"93050400",
		16#1f50# => X"13050900",
		16#1f51# => X"eff09fcd",
		16#1f52# => X"2320a400",
		16#1f53# => X"23200500",
		16#1f54# => X"13040500",
		16#1f55# => X"6ff09ffa",
		16#1f56# => X"8320c101",
		16#1f57# => X"03248101",
		16#1f58# => X"13850900",
		16#1f59# => X"83244101",
		16#1f5a# => X"03290101",
		16#1f5b# => X"8329c100",
		16#1f5c# => X"032a8100",
		16#1f5d# => X"13010102",
		16#1f5e# => X"67800000",
		16#1f5f# => X"130101fd",
		16#1f60# => X"23229102",
		16#1f61# => X"93840500",
		16#1f62# => X"232e3101",
		16#1f63# => X"83a90401",
		16#1f64# => X"23248102",
		16#1f65# => X"83a54500",
		16#1f66# => X"13545640",
		16#1f67# => X"83a78400",
		16#1f68# => X"b3093401",
		16#1f69# => X"23202103",
		16#1f6a# => X"232a5101",
		16#1f6b# => X"23261102",
		16#1f6c# => X"232c4101",
		16#1f6d# => X"930a0500",
		16#1f6e# => X"13891900",
		16#1f6f# => X"63c6270d",
		16#1f70# => X"13850a00",
		16#1f71# => X"2326c100",
		16#1f72# => X"eff08fff",
		16#1f73# => X"0326c100",
		16#1f74# => X"93074501",
		16#1f75# => X"130a0500",
		16#1f76# => X"93860700",
		16#1f77# => X"13070000",
		16#1f78# => X"93864600",
		16#1f79# => X"6348870a",
		16#1f7a# => X"63540400",
		16#1f7b# => X"13040000",
		16#1f7c# => X"83a60401",
		16#1f7d# => X"13142400",
		16#1f7e# => X"33878700",
		16#1f7f# => X"93962600",
		16#1f80# => X"93874401",
		16#1f81# => X"1376f601",
		16#1f82# => X"b386d700",
		16#1f83# => X"630e0608",
		16#1f84# => X"13080002",
		16#1f85# => X"3308c840",
		16#1f86# => X"93050000",
		16#1f87# => X"03a50700",
		16#1f88# => X"93084700",
		16#1f89# => X"93874700",
		16#1f8a# => X"3315c500",
		16#1f8b# => X"b365b500",
		16#1f8c# => X"23aeb8fe",
		16#1f8d# => X"83a5c7ff",
		16#1f8e# => X"b3d50501",
		16#1f8f# => X"63e2d706",
		16#1f90# => X"2322b700",
		16#1f91# => X"63840500",
		16#1f92# => X"13892900",
		16#1f93# => X"1309f9ff",
		16#1f94# => X"23282a01",
		16#1f95# => X"13850a00",
		16#1f96# => X"93850400",
		16#1f97# => X"eff0df80",
		16#1f98# => X"8320c102",
		16#1f99# => X"03248102",
		16#1f9a# => X"13050a00",
		16#1f9b# => X"83244102",
		16#1f9c# => X"03290102",
		16#1f9d# => X"8329c101",
		16#1f9e# => X"032a8101",
		16#1f9f# => X"832a4101",
		16#1fa0# => X"13010103",
		16#1fa1# => X"67800000",
		16#1fa2# => X"93851500",
		16#1fa3# => X"93971700",
		16#1fa4# => X"6ff0dff2",
		16#1fa5# => X"23ae06fe",
		16#1fa6# => X"13071700",
		16#1fa7# => X"6ff05ff4",
		16#1fa8# => X"13870800",
		16#1fa9# => X"6ff09ff7",
		16#1faa# => X"93874700",
		16#1fab# => X"03a6c7ff",
		16#1fac# => X"13074700",
		16#1fad# => X"232ec7fe",
		16#1fae# => X"e3e8d7fe",
		16#1faf# => X"6ff01ff9",
		16#1fb0# => X"83270501",
		16#1fb1# => X"03a70501",
		16#1fb2# => X"b387e740",
		16#1fb3# => X"639c0702",
		16#1fb4# => X"13172700",
		16#1fb5# => X"13054501",
		16#1fb6# => X"93854501",
		16#1fb7# => X"b306e500",
		16#1fb8# => X"b385e500",
		16#1fb9# => X"9386c6ff",
		16#1fba# => X"9385c5ff",
		16#1fbb# => X"03a60600",
		16#1fbc# => X"03a70500",
		16#1fbd# => X"630ce600",
		16#1fbe# => X"9307f0ff",
		16#1fbf# => X"6364e600",
		16#1fc0# => X"93071000",
		16#1fc1# => X"13850700",
		16#1fc2# => X"67800000",
		16#1fc3# => X"e36cd5fc",
		16#1fc4# => X"6ff05fff",
		16#1fc5# => X"130101fe",
		16#1fc6# => X"232a9100",
		16#1fc7# => X"93840500",
		16#1fc8# => X"23263101",
		16#1fc9# => X"93050600",
		16#1fca# => X"93090500",
		16#1fcb# => X"13850400",
		16#1fcc# => X"232c8100",
		16#1fcd# => X"232e1100",
		16#1fce# => X"23282101",
		16#1fcf# => X"13040600",
		16#1fd0# => X"eff01ff8",
		16#1fd1# => X"631c0502",
		16#1fd2# => X"93050000",
		16#1fd3# => X"13850900",
		16#1fd4# => X"eff00fe7",
		16#1fd5# => X"93071000",
		16#1fd6# => X"2328f500",
		16#1fd7# => X"232a0500",
		16#1fd8# => X"8320c101",
		16#1fd9# => X"03248101",
		16#1fda# => X"83244101",
		16#1fdb# => X"03290101",
		16#1fdc# => X"8329c100",
		16#1fdd# => X"13010102",
		16#1fde# => X"67800000",
		16#1fdf# => X"13091000",
		16#1fe0# => X"634a0500",
		16#1fe1# => X"93070400",
		16#1fe2# => X"13090000",
		16#1fe3# => X"13840400",
		16#1fe4# => X"93840700",
		16#1fe5# => X"83254400",
		16#1fe6# => X"13850900",
		16#1fe7# => X"eff04fe2",
		16#1fe8# => X"03230401",
		16#1fe9# => X"83a80401",
		16#1fea# => X"13064401",
		16#1feb# => X"131e2300",
		16#1fec# => X"13884401",
		16#1fed# => X"93982800",
		16#1fee# => X"b70e0100",
		16#1fef# => X"23262501",
		16#1ff0# => X"330ec601",
		16#1ff1# => X"b3081801",
		16#1ff2# => X"93064501",
		16#1ff3# => X"130f0000",
		16#1ff4# => X"938efeff",
		16#1ff5# => X"03270600",
		16#1ff6# => X"832f0800",
		16#1ff7# => X"93864600",
		16#1ff8# => X"b375d701",
		16#1ff9# => X"b3f7df01",
		16#1ffa# => X"b385e501",
		16#1ffb# => X"b385f540",
		16#1ffc# => X"93df0f01",
		16#1ffd# => X"93570701",
		16#1ffe# => X"b387f741",
		16#1fff# => X"13d70541",
		16#2000# => X"b387e700",
		16#2001# => X"13df0741",
		16#2002# => X"b3f5d501",
		16#2003# => X"93970701",
		16#2004# => X"b3e7b700",
		16#2005# => X"13084800",
		16#2006# => X"23aef6fe",
		16#2007# => X"13064600",
		16#2008# => X"e36a18fb",
		16#2009# => X"b7050100",
		16#200a# => X"9385f5ff",
		16#200b# => X"636cc601",
		16#200c# => X"9386c6ff",
		16#200d# => X"83a70600",
		16#200e# => X"63820704",
		16#200f# => X"23286500",
		16#2010# => X"6ff01ff2",
		16#2011# => X"83270600",
		16#2012# => X"93864600",
		16#2013# => X"13064600",
		16#2014# => X"33f7b700",
		16#2015# => X"3307e701",
		16#2016# => X"13580741",
		16#2017# => X"93d70701",
		16#2018# => X"b3870701",
		16#2019# => X"13df0741",
		16#201a# => X"3377b700",
		16#201b# => X"93970701",
		16#201c# => X"b3e7e700",
		16#201d# => X"23aef6fe",
		16#201e# => X"6ff05ffb",
		16#201f# => X"1303f3ff",
		16#2020# => X"6ff01ffb",
		16#2021# => X"b707f07f",
		16#2022# => X"b3f5b700",
		16#2023# => X"b707c0fc",
		16#2024# => X"b385f500",
		16#2025# => X"6358b000",
		16#2026# => X"93070000",
		16#2027# => X"13850700",
		16#2028# => X"67800000",
		16#2029# => X"b305b040",
		16#202a# => X"93d74541",
		16#202b# => X"13073001",
		16#202c# => X"6348f700",
		16#202d# => X"b7050800",
		16#202e# => X"b3d5f540",
		16#202f# => X"6ff0dffd",
		16#2030# => X"9387c7fe",
		16#2031# => X"9306e001",
		16#2032# => X"93050000",
		16#2033# => X"13071000",
		16#2034# => X"63c6f600",
		16#2035# => X"93c7f7ff",
		16#2036# => X"3317f700",
		16#2037# => X"93070700",
		16#2038# => X"6ff0dffb",
		16#2039# => X"130101fd",
		16#203a# => X"23229102",
		16#203b# => X"83240501",
		16#203c# => X"232e3101",
		16#203d# => X"93094501",
		16#203e# => X"93942400",
		16#203f# => X"b3849900",
		16#2040# => X"23248102",
		16#2041# => X"03a4c4ff",
		16#2042# => X"23202103",
		16#2043# => X"2326b100",
		16#2044# => X"13050400",
		16#2045# => X"23261102",
		16#2046# => X"eff0cffa",
		16#2047# => X"8325c100",
		16#2048# => X"93070002",
		16#2049# => X"b387a740",
		16#204a# => X"23a0f500",
		16#204b# => X"9307a000",
		16#204c# => X"1389c4ff",
		16#204d# => X"63cca704",
		16#204e# => X"9307b000",
		16#204f# => X"b387a740",
		16#2050# => X"3707f03f",
		16#2051# => X"b356f400",
		16#2052# => X"b3e6e600",
		16#2053# => X"13070000",
		16#2054# => X"63f42901",
		16#2055# => X"03a784ff",
		16#2056# => X"13055501",
		16#2057# => X"3315a400",
		16#2058# => X"b357f700",
		16#2059# => X"b367f500",
		16#205a# => X"8320c102",
		16#205b# => X"03248102",
		16#205c# => X"83244102",
		16#205d# => X"03290102",
		16#205e# => X"8329c101",
		16#205f# => X"13850700",
		16#2060# => X"93850600",
		16#2061# => X"13010103",
		16#2062# => X"67800000",
		16#2063# => X"93070000",
		16#2064# => X"63f62901",
		16#2065# => X"83a784ff",
		16#2066# => X"138984ff",
		16#2067# => X"130555ff",
		16#2068# => X"630e0502",
		16#2069# => X"13070002",
		16#206a# => X"3306a740",
		16#206b# => X"3314a400",
		16#206c# => X"3707f03f",
		16#206d# => X"3364e400",
		16#206e# => X"b3d6c700",
		16#206f# => X"b366d400",
		16#2070# => X"13070000",
		16#2071# => X"63f42901",
		16#2072# => X"0327c9ff",
		16#2073# => X"b397a700",
		16#2074# => X"3357c700",
		16#2075# => X"b3e7e700",
		16#2076# => X"6ff01ff9",
		16#2077# => X"b706f03f",
		16#2078# => X"b366d400",
		16#2079# => X"6ff05ff8",
		16#207a# => X"130101fd",
		16#207b# => X"23248102",
		16#207c# => X"13840500",
		16#207d# => X"93051000",
		16#207e# => X"23229102",
		16#207f# => X"23202103",
		16#2080# => X"93040600",
		16#2081# => X"232e3101",
		16#2082# => X"232c4101",
		16#2083# => X"13090700",
		16#2084# => X"23261102",
		16#2085# => X"138a0600",
		16#2086# => X"eff08fba",
		16#2087# => X"37071000",
		16#2088# => X"9307f7ff",
		16#2089# => X"b3f79700",
		16#208a# => X"93d44401",
		16#208b# => X"93f4f47f",
		16#208c# => X"93090500",
		16#208d# => X"639a0408",
		16#208e# => X"2326f100",
		16#208f# => X"630e0408",
		16#2090# => X"13058100",
		16#2091# => X"23248100",
		16#2092# => X"eff00fef",
		16#2093# => X"83268100",
		16#2094# => X"63000508",
		16#2095# => X"0327c100",
		16#2096# => X"93070002",
		16#2097# => X"b387a740",
		16#2098# => X"b317f700",
		16#2099# => X"b3e7d700",
		16#209a# => X"3357a700",
		16#209b# => X"23aaf900",
		16#209c# => X"2326e100",
		16#209d# => X"0324c100",
		16#209e# => X"23ac8900",
		16#209f# => X"33348000",
		16#20a0# => X"13041400",
		16#20a1# => X"23a88900",
		16#20a2# => X"638a0406",
		16#20a3# => X"9384d4bc",
		16#20a4# => X"b384a400",
		16#20a5# => X"93075003",
		16#20a6# => X"23209a00",
		16#20a7# => X"3385a740",
		16#20a8# => X"2320a900",
		16#20a9# => X"8320c102",
		16#20aa# => X"03248102",
		16#20ab# => X"13850900",
		16#20ac# => X"83244102",
		16#20ad# => X"03290102",
		16#20ae# => X"8329c101",
		16#20af# => X"032a8101",
		16#20b0# => X"13010103",
		16#20b1# => X"67800000",
		16#20b2# => X"b3e7e700",
		16#20b3# => X"6ff0dff6",
		16#20b4# => X"23aad900",
		16#20b5# => X"6ff01ffa",
		16#20b6# => X"1305c100",
		16#20b7# => X"eff0cfe5",
		16#20b8# => X"8327c100",
		16#20b9# => X"13050502",
		16#20ba# => X"13041000",
		16#20bb# => X"23aaf900",
		16#20bc# => X"93071000",
		16#20bd# => X"23a8f900",
		16#20be# => X"6ff01ff9",
		16#20bf# => X"93172400",
		16#20c0# => X"1305e5bc",
		16#20c1# => X"b387f900",
		16#20c2# => X"2320aa00",
		16#20c3# => X"03a50701",
		16#20c4# => X"13145400",
		16#20c5# => X"eff00fdb",
		16#20c6# => X"3304a440",
		16#20c7# => X"23208900",
		16#20c8# => X"6ff05ff8",
		16#20c9# => X"130101fd",
		16#20ca# => X"232c4101",
		16#20cb# => X"138a0500",
		16#20cc# => X"93058100",
		16#20cd# => X"23261102",
		16#20ce# => X"23248102",
		16#20cf# => X"23229102",
		16#20d0# => X"232e3101",
		16#20d1# => X"232a5101",
		16#20d2# => X"23286101",
		16#20d3# => X"23202103",
		16#20d4# => X"130b0500",
		16#20d5# => X"eff01fd9",
		16#20d6# => X"13040500",
		16#20d7# => X"93890500",
		16#20d8# => X"93840500",
		16#20d9# => X"13050a00",
		16#20da# => X"9305c100",
		16#20db# => X"eff09fd7",
		16#20dc# => X"930a0500",
		16#20dd# => X"83270b01",
		16#20de# => X"03250a01",
		16#20df# => X"0327c100",
		16#20e0# => X"b387a740",
		16#20e1# => X"03258100",
		16#20e2# => X"93975700",
		16#20e3# => X"3305e540",
		16#20e4# => X"3385a700",
		16#20e5# => X"6358a004",
		16#20e6# => X"13154501",
		16#20e7# => X"93860500",
		16#20e8# => X"b3043501",
		16#20e9# => X"93870600",
		16#20ea# => X"13860a00",
		16#20eb# => X"13050400",
		16#20ec# => X"93850400",
		16#20ed# => X"93860700",
		16#20ee# => X"ef509060",
		16#20ef# => X"8320c102",
		16#20f0# => X"03248102",
		16#20f1# => X"83244102",
		16#20f2# => X"03290102",
		16#20f3# => X"8329c101",
		16#20f4# => X"032a8101",
		16#20f5# => X"832a4101",
		16#20f6# => X"032b0101",
		16#20f7# => X"13010103",
		16#20f8# => X"67800000",
		16#20f9# => X"13890500",
		16#20fa# => X"b705f0ff",
		16#20fb# => X"efa04024",
		16#20fc# => X"b3062501",
		16#20fd# => X"6ff01ffb",
		16#20fe# => X"130101ff",
		16#20ff# => X"23248100",
		16#2100# => X"23261100",
		16#2101# => X"23222101",
		16#2102# => X"23203101",
		16#2103# => X"93077001",
		16#2104# => X"13040500",
		16#2105# => X"63caa702",
		16#2106# => X"b7470110",
		16#2107# => X"13143500",
		16#2108# => X"938787f3",
		16#2109# => X"33848700",
		16#210a# => X"03250401",
		16#210b# => X"83254401",
		16#210c# => X"8320c100",
		16#210d# => X"03248100",
		16#210e# => X"03294100",
		16#210f# => X"83290100",
		16#2110# => X"13010101",
		16#2111# => X"67800000",
		16#2112# => X"b7570110",
		16#2113# => X"03a58721",
		16#2114# => X"83a5c721",
		16#2115# => X"b7570110",
		16#2116# => X"03a90722",
		16#2117# => X"83a94722",
		16#2118# => X"13060900",
		16#2119# => X"93860900",
		16#211a# => X"1304f4ff",
		16#211b# => X"ef600056",
		16#211c# => X"e31804fe",
		16#211d# => X"6ff0dffb",
		16#211e# => X"9387f5ff",
		16#211f# => X"03270601",
		16#2120# => X"93d75740",
		16#2121# => X"93871700",
		16#2122# => X"93972700",
		16#2123# => X"93064601",
		16#2124# => X"13172700",
		16#2125# => X"b307f500",
		16#2126# => X"3387e600",
		16#2127# => X"63e6e600",
		16#2128# => X"636ef500",
		16#2129# => X"67800000",
		16#212a# => X"93864600",
		16#212b# => X"03a6c6ff",
		16#212c# => X"13054500",
		16#212d# => X"232ec5fe",
		16#212e# => X"6ff05ffe",
		16#212f# => X"13054500",
		16#2130# => X"232e05fe",
		16#2131# => X"6ff0dffd",
		16#2132# => X"83260501",
		16#2133# => X"93d75540",
		16#2134# => X"13074501",
		16#2135# => X"63c0f604",
		16#2136# => X"63d4d702",
		16#2137# => X"93f5f501",
		16#2138# => X"63800502",
		16#2139# => X"93962700",
		16#213a# => X"b306d700",
		16#213b# => X"03a60600",
		16#213c# => X"13051000",
		16#213d# => X"b356b600",
		16#213e# => X"b395b600",
		16#213f# => X"6318b602",
		16#2140# => X"93972700",
		16#2141# => X"b307f700",
		16#2142# => X"636af700",
		16#2143# => X"13050000",
		16#2144# => X"67800000",
		16#2145# => X"93870600",
		16#2146# => X"6ff09ffe",
		16#2147# => X"9387c7ff",
		16#2148# => X"83a60700",
		16#2149# => X"e38206fe",
		16#214a# => X"13051000",
		16#214b# => X"67800000",
		16#214c# => X"130101fc",
		16#214d# => X"232c8102",
		16#214e# => X"232e1102",
		16#214f# => X"13840500",
		16#2150# => X"232a9102",
		16#2151# => X"23282103",
		16#2152# => X"23263103",
		16#2153# => X"23244103",
		16#2154# => X"23225103",
		16#2155# => X"23206103",
		16#2156# => X"232e7101",
		16#2157# => X"232c8101",
		16#2158# => X"93050600",
		16#2159# => X"631a0402",
		16#215a# => X"03248103",
		16#215b# => X"8320c103",
		16#215c# => X"83244103",
		16#215d# => X"03290103",
		16#215e# => X"8329c102",
		16#215f# => X"032a8102",
		16#2160# => X"832a4102",
		16#2161# => X"032b0102",
		16#2162# => X"832bc101",
		16#2163# => X"032c8101",
		16#2164# => X"13010104",
		16#2165# => X"6fe04ff2",
		16#2166# => X"930a0500",
		16#2167# => X"2326c100",
		16#2168# => X"eff08f81",
		16#2169# => X"8325c100",
		16#216a# => X"8326c4ff",
		16#216b# => X"93076001",
		16#216c# => X"9389b500",
		16#216d# => X"930b84ff",
		16#216e# => X"13f9c6ff",
		16#216f# => X"63f63705",
		16#2170# => X"13fb89ff",
		16#2171# => X"63540b04",
		16#2172# => X"9307c000",
		16#2173# => X"23a0fa00",
		16#2174# => X"130a0000",
		16#2175# => X"8320c103",
		16#2176# => X"03248103",
		16#2177# => X"13050a00",
		16#2178# => X"83244103",
		16#2179# => X"03290103",
		16#217a# => X"8329c102",
		16#217b# => X"032a8102",
		16#217c# => X"832a4102",
		16#217d# => X"032b0102",
		16#217e# => X"832bc101",
		16#217f# => X"032c8101",
		16#2180# => X"13010104",
		16#2181# => X"67800000",
		16#2182# => X"130b0001",
		16#2183# => X"e36ebbfa",
		16#2184# => X"635c6945",
		16#2185# => X"375c0110",
		16#2186# => X"1307cce0",
		16#2187# => X"03268700",
		16#2188# => X"b3872b01",
		16#2189# => X"03a74700",
		16#218a# => X"130ccce0",
		16#218b# => X"630cf600",
		16#218c# => X"1375e7ff",
		16#218d# => X"3385a700",
		16#218e# => X"03254500",
		16#218f# => X"13751500",
		16#2190# => X"631a050a",
		16#2191# => X"1377c7ff",
		16#2192# => X"b309e900",
		16#2193# => X"6310f604",
		16#2194# => X"13050b01",
		16#2195# => X"63c4a90a",
		16#2196# => X"b38b6b01",
		16#2197# => X"b3896941",
		16#2198# => X"23247c01",
		16#2199# => X"93e91900",
		16#219a# => X"23a23b01",
		16#219b# => X"8329c4ff",
		16#219c# => X"13850a00",
		16#219d# => X"130a0400",
		16#219e# => X"93f91900",
		16#219f# => X"b3e96901",
		16#21a0# => X"232e34ff",
		16#21a1# => X"efe09ff3",
		16#21a2# => X"6ff0dff4",
		16#21a3# => X"63c86907",
		16#21a4# => X"03a7c700",
		16#21a5# => X"83a78700",
		16#21a6# => X"23a6e700",
		16#21a7# => X"2324f700",
		16#21a8# => X"03a74b00",
		16#21a9# => X"b3866941",
		16#21aa# => X"1306f000",
		16#21ab# => X"13771700",
		16#21ac# => X"b3873b01",
		16#21ad# => X"637ed63a",
		16#21ae# => X"b369eb00",
		16#21af# => X"23a23b01",
		16#21b0# => X"b3856b01",
		16#21b1# => X"93e61600",
		16#21b2# => X"23a2d500",
		16#21b3# => X"03a74700",
		16#21b4# => X"93858500",
		16#21b5# => X"13850a00",
		16#21b6# => X"13671700",
		16#21b7# => X"23a2e700",
		16#21b8# => X"efb0dfab",
		16#21b9# => X"13850a00",
		16#21ba# => X"efe05fed",
		16#21bb# => X"138a8b00",
		16#21bc# => X"6ff05fee",
		16#21bd# => X"13070000",
		16#21be# => X"93070000",
		16#21bf# => X"93f61600",
		16#21c0# => X"63920628",
		16#21c1# => X"832484ff",
		16#21c2# => X"b3849b40",
		16#21c3# => X"03aa4400",
		16#21c4# => X"137acaff",
		16#21c5# => X"330a2a01",
		16#21c6# => X"638c071a",
		16#21c7# => X"b3094701",
		16#21c8# => X"6316f60e",
		16#21c9# => X"93070b01",
		16#21ca# => X"63c4f91a",
		16#21cb# => X"03a78400",
		16#21cc# => X"83a7c400",
		16#21cd# => X"1306c9ff",
		16#21ce# => X"138a8400",
		16#21cf# => X"2326f700",
		16#21d0# => X"23a4e700",
		16#21d1# => X"13074002",
		16#21d2# => X"636ac70a",
		16#21d3# => X"93063001",
		16#21d4# => X"93070a00",
		16#21d5# => X"63f2c602",
		16#21d6# => X"83270400",
		16#21d7# => X"23a4f400",
		16#21d8# => X"83274400",
		16#21d9# => X"23a6f400",
		16#21da# => X"9307b001",
		16#21db# => X"63eac704",
		16#21dc# => X"13048400",
		16#21dd# => X"93870401",
		16#21de# => X"03270400",
		16#21df# => X"23a0e700",
		16#21e0# => X"03274400",
		16#21e1# => X"23a2e700",
		16#21e2# => X"03278400",
		16#21e3# => X"23a4e700",
		16#21e4# => X"b3876401",
		16#21e5# => X"b3896941",
		16#21e6# => X"2324fc00",
		16#21e7# => X"93e91900",
		16#21e8# => X"23a23701",
		16#21e9# => X"83a74400",
		16#21ea# => X"93f71700",
		16#21eb# => X"b3e96701",
		16#21ec# => X"23a23401",
		16#21ed# => X"13850a00",
		16#21ee# => X"efe05fe0",
		16#21ef# => X"6ff09fe1",
		16#21f0# => X"83278400",
		16#21f1# => X"23a8f400",
		16#21f2# => X"8327c400",
		16#21f3# => X"23aaf400",
		16#21f4# => X"6308e600",
		16#21f5# => X"13040401",
		16#21f6# => X"93878401",
		16#21f7# => X"6ff0dff9",
		16#21f8# => X"83270401",
		16#21f9# => X"13048401",
		16#21fa# => X"23acf400",
		16#21fb# => X"0327c4ff",
		16#21fc# => X"93870402",
		16#21fd# => X"23aee400",
		16#21fe# => X"6ff01ff8",
		16#21ff# => X"93050400",
		16#2200# => X"13050a00",
		16#2201# => X"efe05fc8",
		16#2202# => X"6ff09ff8",
		16#2203# => X"63c2690d",
		16#2204# => X"03a7c700",
		16#2205# => X"83a78700",
		16#2206# => X"1306c9ff",
		16#2207# => X"13858400",
		16#2208# => X"23a6e700",
		16#2209# => X"2324f700",
		16#220a# => X"03a78400",
		16#220b# => X"83a7c400",
		16#220c# => X"2326f700",
		16#220d# => X"23a4e700",
		16#220e# => X"93074002",
		16#220f# => X"63e4c708",
		16#2210# => X"13073001",
		16#2211# => X"6372c702",
		16#2212# => X"03270400",
		16#2213# => X"23a4e400",
		16#2214# => X"03274400",
		16#2215# => X"23a6e400",
		16#2216# => X"1307b001",
		16#2217# => X"6366c702",
		16#2218# => X"13048400",
		16#2219# => X"13850401",
		16#221a# => X"83270400",
		16#221b# => X"2320f500",
		16#221c# => X"83274400",
		16#221d# => X"2322f500",
		16#221e# => X"83278400",
		16#221f# => X"2324f500",
		16#2220# => X"938b0400",
		16#2221# => X"6ff0dfe1",
		16#2222# => X"03278400",
		16#2223# => X"23a8e400",
		16#2224# => X"0327c400",
		16#2225# => X"23aae400",
		16#2226# => X"6308f600",
		16#2227# => X"13040401",
		16#2228# => X"13858401",
		16#2229# => X"6ff05ffc",
		16#222a# => X"83270401",
		16#222b# => X"13850402",
		16#222c# => X"13048401",
		16#222d# => X"23acf400",
		16#222e# => X"8327c4ff",
		16#222f# => X"23aef400",
		16#2230# => X"6ff09ffa",
		16#2231# => X"93050400",
		16#2232# => X"efe01fbc",
		16#2233# => X"6ff05ffb",
		16#2234# => X"634a6a0b",
		16#2235# => X"83a7c400",
		16#2236# => X"03a78400",
		16#2237# => X"1306c9ff",
		16#2238# => X"13858400",
		16#2239# => X"2326f700",
		16#223a# => X"23a4e700",
		16#223b# => X"93074002",
		16#223c# => X"63e4c708",
		16#223d# => X"13073001",
		16#223e# => X"6372c702",
		16#223f# => X"03270400",
		16#2240# => X"23a4e400",
		16#2241# => X"03274400",
		16#2242# => X"23a6e400",
		16#2243# => X"1307b001",
		16#2244# => X"6366c702",
		16#2245# => X"13048400",
		16#2246# => X"13850401",
		16#2247# => X"83270400",
		16#2248# => X"2320f500",
		16#2249# => X"83274400",
		16#224a# => X"2322f500",
		16#224b# => X"83278400",
		16#224c# => X"2324f500",
		16#224d# => X"93090a00",
		16#224e# => X"6ff09ff4",
		16#224f# => X"03278400",
		16#2250# => X"23a8e400",
		16#2251# => X"0327c400",
		16#2252# => X"23aae400",
		16#2253# => X"6308f600",
		16#2254# => X"13040401",
		16#2255# => X"13858401",
		16#2256# => X"6ff05ffc",
		16#2257# => X"83270401",
		16#2258# => X"13850402",
		16#2259# => X"13048401",
		16#225a# => X"23acf400",
		16#225b# => X"8327c4ff",
		16#225c# => X"23aef400",
		16#225d# => X"6ff09ffa",
		16#225e# => X"93050400",
		16#225f# => X"efe0dfb0",
		16#2260# => X"6ff05ffb",
		16#2261# => X"13850a00",
		16#2262# => X"efe00fb3",
		16#2263# => X"130a0500",
		16#2264# => X"e30205e2",
		16#2265# => X"8327c4ff",
		16#2266# => X"130785ff",
		16#2267# => X"93f7e7ff",
		16#2268# => X"b387fb00",
		16#2269# => X"639ae700",
		16#226a# => X"8329c5ff",
		16#226b# => X"93f9c9ff",
		16#226c# => X"b3892901",
		16#226d# => X"6ff0dfce",
		16#226e# => X"1306c9ff",
		16#226f# => X"93074002",
		16#2270# => X"63eec708",
		16#2271# => X"13073001",
		16#2272# => X"6374c708",
		16#2273# => X"03270400",
		16#2274# => X"2320e500",
		16#2275# => X"03274400",
		16#2276# => X"2322e500",
		16#2277# => X"1307b001",
		16#2278# => X"636ac702",
		16#2279# => X"13078400",
		16#227a# => X"93078500",
		16#227b# => X"83260700",
		16#227c# => X"23a0d700",
		16#227d# => X"83264700",
		16#227e# => X"23a2d700",
		16#227f# => X"03278700",
		16#2280# => X"23a4e700",
		16#2281# => X"93050400",
		16#2282# => X"13850a00",
		16#2283# => X"efb00ff9",
		16#2284# => X"6ff05fda",
		16#2285# => X"03278400",
		16#2286# => X"2324e500",
		16#2287# => X"0327c400",
		16#2288# => X"2326e500",
		16#2289# => X"6308f600",
		16#228a# => X"13070401",
		16#228b# => X"93070501",
		16#228c# => X"6ff0dffb",
		16#228d# => X"83270401",
		16#228e# => X"13078401",
		16#228f# => X"2328f500",
		16#2290# => X"83264401",
		16#2291# => X"93078501",
		16#2292# => X"232ad500",
		16#2293# => X"6ff01ffa",
		16#2294# => X"93070500",
		16#2295# => X"13070400",
		16#2296# => X"6ff05ff9",
		16#2297# => X"93050400",
		16#2298# => X"efe09fa2",
		16#2299# => X"6ff01ffa",
		16#229a# => X"93090900",
		16#229b# => X"6ff05fc3",
		16#229c# => X"b3e9e900",
		16#229d# => X"23a23b01",
		16#229e# => X"03a74700",
		16#229f# => X"13671700",
		16#22a0# => X"23a2e700",
		16#22a1# => X"6ff01fc6",
		16#22a2# => X"130101ff",
		16#22a3# => X"23248100",
		16#22a4# => X"23229100",
		16#22a5# => X"37840110",
		16#22a6# => X"93040500",
		16#22a7# => X"13850500",
		16#22a8# => X"23261100",
		16#22a9# => X"232204aa",
		16#22aa# => X"ef40d027",
		16#22ab# => X"9307f0ff",
		16#22ac# => X"6318f500",
		16#22ad# => X"832744aa",
		16#22ae# => X"63840700",
		16#22af# => X"23a0f400",
		16#22b0# => X"8320c100",
		16#22b1# => X"03248100",
		16#22b2# => X"83244100",
		16#22b3# => X"13010101",
		16#22b4# => X"67800000",
		16#22b5# => X"130101ff",
		16#22b6# => X"23229100",
		16#22b7# => X"b7040080",
		16#22b8# => X"23248100",
		16#22b9# => X"23261100",
		16#22ba# => X"93c4f4ff",
		16#22bb# => X"33f7b400",
		16#22bc# => X"23200600",
		16#22bd# => X"3708f07f",
		16#22be# => X"93060500",
		16#22bf# => X"93870500",
		16#22c0# => X"13040600",
		16#22c1# => X"63520707",
		16#22c2# => X"3368a700",
		16#22c3# => X"630e0804",
		16#22c4# => X"b7071000",
		16#22c5# => X"13860500",
		16#22c6# => X"6354f702",
		16#22c7# => X"b7570110",
		16#22c8# => X"03a68722",
		16#22c9# => X"83a6c722",
		16#22ca# => X"ef50506a",
		16#22cb# => X"9307a0fc",
		16#22cc# => X"93060500",
		16#22cd# => X"13860500",
		16#22ce# => X"33f7b400",
		16#22cf# => X"2320f400",
		16#22d0# => X"83270400",
		16#22d1# => X"13574741",
		16#22d2# => X"130727c0",
		16#22d3# => X"3387e700",
		16#22d4# => X"b7071080",
		16#22d5# => X"9387f7ff",
		16#22d6# => X"3376f600",
		16#22d7# => X"b707e03f",
		16#22d8# => X"2320e400",
		16#22d9# => X"b367f600",
		16#22da# => X"8320c100",
		16#22db# => X"03248100",
		16#22dc# => X"83244100",
		16#22dd# => X"13850600",
		16#22de# => X"93850700",
		16#22df# => X"13010101",
		16#22e0# => X"67800000",
		16#22e1# => X"130101f6",
		16#22e2# => X"232af108",
		16#22e3# => X"b7070080",
		16#22e4# => X"93c7f7ff",
		16#22e5# => X"232ef100",
		16#22e6# => X"2328f100",
		16#22e7# => X"b707ffff",
		16#22e8# => X"2326d108",
		16#22e9# => X"2324b100",
		16#22ea# => X"232cb100",
		16#22eb# => X"93878720",
		16#22ec# => X"9306c108",
		16#22ed# => X"93058100",
		16#22ee# => X"232e1106",
		16#22ef# => X"232af100",
		16#22f0# => X"2328e108",
		16#22f1# => X"232c0109",
		16#22f2# => X"232e1109",
		16#22f3# => X"2322d100",
		16#22f4# => X"ef008022",
		16#22f5# => X"83278100",
		16#22f6# => X"23800700",
		16#22f7# => X"8320c107",
		16#22f8# => X"1301010a",
		16#22f9# => X"67800000",
		16#22fa# => X"130101f6",
		16#22fb# => X"232af108",
		16#22fc# => X"b7070080",
		16#22fd# => X"93c7f7ff",
		16#22fe# => X"232ef100",
		16#22ff# => X"2328f100",
		16#2300# => X"b707ffff",
		16#2301# => X"93878720",
		16#2302# => X"232af100",
		16#2303# => X"2324a100",
		16#2304# => X"232ca100",
		16#2305# => X"03a5c181",
		16#2306# => X"2324c108",
		16#2307# => X"2326d108",
		16#2308# => X"13860500",
		16#2309# => X"93068108",
		16#230a# => X"93058100",
		16#230b# => X"232e1106",
		16#230c# => X"2328e108",
		16#230d# => X"232c0109",
		16#230e# => X"232e1109",
		16#230f# => X"2322d100",
		16#2310# => X"ef00801b",
		16#2311# => X"83278100",
		16#2312# => X"23800700",
		16#2313# => X"8320c107",
		16#2314# => X"1301010a",
		16#2315# => X"67800000",
		16#2316# => X"130101ff",
		16#2317# => X"23248100",
		16#2318# => X"13840500",
		16#2319# => X"8395e500",
		16#231a# => X"23261100",
		16#231b# => X"ef304043",
		16#231c# => X"63400502",
		16#231d# => X"83270405",
		16#231e# => X"b387a700",
		16#231f# => X"2328f404",
		16#2320# => X"8320c100",
		16#2321# => X"03248100",
		16#2322# => X"13010101",
		16#2323# => X"67800000",
		16#2324# => X"8357c400",
		16#2325# => X"37f7ffff",
		16#2326# => X"1307f7ff",
		16#2327# => X"b3f7e700",
		16#2328# => X"2316f400",
		16#2329# => X"6ff0dffd",
		16#232a# => X"13050000",
		16#232b# => X"67800000",
		16#232c# => X"83d7c500",
		16#232d# => X"130101fe",
		16#232e# => X"232c8100",
		16#232f# => X"232a9100",
		16#2330# => X"23282101",
		16#2331# => X"23263101",
		16#2332# => X"232e1100",
		16#2333# => X"93f70710",
		16#2334# => X"93040500",
		16#2335# => X"13840500",
		16#2336# => X"13090600",
		16#2337# => X"93890600",
		16#2338# => X"638a0700",
		16#2339# => X"8395e500",
		16#233a# => X"93062000",
		16#233b# => X"13060000",
		16#233c# => X"ef30c035",
		16#233d# => X"8357c400",
		16#233e# => X"37f7ffff",
		16#233f# => X"1307f7ff",
		16#2340# => X"b3f7e700",
		16#2341# => X"2316f400",
		16#2342# => X"8315e400",
		16#2343# => X"03248101",
		16#2344# => X"8320c101",
		16#2345# => X"93860900",
		16#2346# => X"13060900",
		16#2347# => X"8329c100",
		16#2348# => X"03290101",
		16#2349# => X"13850400",
		16#234a# => X"83244101",
		16#234b# => X"13010102",
		16#234c# => X"6f20506b",
		16#234d# => X"130101ff",
		16#234e# => X"23248100",
		16#234f# => X"13840500",
		16#2350# => X"8395e500",
		16#2351# => X"23261100",
		16#2352# => X"ef304030",
		16#2353# => X"9307f0ff",
		16#2354# => X"0357c400",
		16#2355# => X"6312f502",
		16#2356# => X"b7f7ffff",
		16#2357# => X"9387f7ff",
		16#2358# => X"b3f7e700",
		16#2359# => X"2316f400",
		16#235a# => X"8320c100",
		16#235b# => X"03248100",
		16#235c# => X"13010101",
		16#235d# => X"67800000",
		16#235e# => X"b7170000",
		16#235f# => X"b367f700",
		16#2360# => X"2316f400",
		16#2361# => X"2328a404",
		16#2362# => X"6ff01ffe",
		16#2363# => X"8395e500",
		16#2364# => X"6f209075",
		16#2365# => X"93070500",
		16#2366# => X"03c70500",
		16#2367# => X"93871700",
		16#2368# => X"93851500",
		16#2369# => X"a38fe7fe",
		16#236a# => X"e31807fe",
		16#236b# => X"67800000",
		16#236c# => X"13070500",
		16#236d# => X"63140600",
		16#236e# => X"67800000",
		16#236f# => X"93851500",
		16#2370# => X"83c6f5ff",
		16#2371# => X"93071700",
		16#2372# => X"1308f6ff",
		16#2373# => X"a38fd7fe",
		16#2374# => X"63980600",
		16#2375# => X"3307c700",
		16#2376# => X"639ae700",
		16#2377# => X"67800000",
		16#2378# => X"13870700",
		16#2379# => X"13060800",
		16#237a# => X"6ff0dffc",
		16#237b# => X"93871700",
		16#237c# => X"a38f07fe",
		16#237d# => X"6ff05ffe",
		16#237e# => X"130101e2",
		16#237f# => X"232e111c",
		16#2380# => X"232a911c",
		16#2381# => X"2328211d",
		16#2382# => X"2326311d",
		16#2383# => X"232c811b",
		16#2384# => X"93890500",
		16#2385# => X"93040600",
		16#2386# => X"138c0600",
		16#2387# => X"232c811c",
		16#2388# => X"2324411d",
		16#2389# => X"2322511d",
		16#238a# => X"2320611d",
		16#238b# => X"232e711b",
		16#238c# => X"232a911b",
		16#238d# => X"2328a11b",
		16#238e# => X"2326b11b",
		16#238f# => X"13090500",
		16#2390# => X"efd01fbf",
		16#2391# => X"83270500",
		16#2392# => X"13850700",
		16#2393# => X"232cf102",
		16#2394# => X"ef805f9c",
		16#2395# => X"83d7c900",
		16#2396# => X"2322a102",
		16#2397# => X"2320010e",
		16#2398# => X"2322010e",
		16#2399# => X"2324010e",
		16#239a# => X"2326010e",
		16#239b# => X"93f70708",
		16#239c# => X"63800704",
		16#239d# => X"83a70901",
		16#239e# => X"639c0702",
		16#239f# => X"93050004",
		16#23a0# => X"13050900",
		16#23a1# => X"efd05fe3",
		16#23a2# => X"23a0a900",
		16#23a3# => X"23a8a900",
		16#23a4# => X"631c0500",
		16#23a5# => X"9307c000",
		16#23a6# => X"2320f900",
		16#23a7# => X"9307f0ff",
		16#23a8# => X"2324f102",
		16#23a9# => X"6f009004",
		16#23aa# => X"93070004",
		16#23ab# => X"23aaf900",
		16#23ac# => X"b7470110",
		16#23ad# => X"93870706",
		16#23ae# => X"2328f104",
		16#23af# => X"b7470110",
		16#23b0# => X"9308c10f",
		16#23b1# => X"9387c71d",
		16#23b2# => X"232a110d",
		16#23b3# => X"232e010c",
		16#23b4# => X"232c010c",
		16#23b5# => X"130a0000",
		16#23b6# => X"138d0800",
		16#23b7# => X"23220104",
		16#23b8# => X"23200104",
		16#23b9# => X"232a0100",
		16#23ba# => X"232a0102",
		16#23bb# => X"232e0102",
		16#23bc# => X"23240102",
		16#23bd# => X"232cf100",
		16#23be# => X"13840400",
		16#23bf# => X"13075002",
		16#23c0# => X"83470400",
		16#23c1# => X"63840700",
		16#23c2# => X"6392e70c",
		16#23c3# => X"b30a9440",
		16#23c4# => X"638a0a04",
		16#23c5# => X"8327c10d",
		16#23c6# => X"23209d00",
		16#23c7# => X"23225d01",
		16#23c8# => X"b3875701",
		16#23c9# => X"232ef10c",
		16#23ca# => X"8327810d",
		16#23cb# => X"13077000",
		16#23cc# => X"130d8d00",
		16#23cd# => X"93871700",
		16#23ce# => X"232cf10c",
		16#23cf# => X"635ef700",
		16#23d0# => X"1306410d",
		16#23d1# => X"93850900",
		16#23d2# => X"13050900",
		16#23d3# => X"ef30402f",
		16#23d4# => X"63180578",
		16#23d5# => X"130dc10f",
		16#23d6# => X"83278102",
		16#23d7# => X"b3875701",
		16#23d8# => X"2324f102",
		16#23d9# => X"83470400",
		16#23da# => X"63940700",
		16#23db# => X"6f10d05c",
		16#23dc# => X"93071400",
		16#23dd# => X"2320f102",
		16#23de# => X"a30b010a",
		16#23df# => X"130bf0ff",
		16#23e0# => X"23260102",
		16#23e1# => X"13040000",
		16#23e2# => X"930a9000",
		16#23e3# => X"930ba005",
		16#23e4# => X"83270102",
		16#23e5# => X"83c70700",
		16#23e6# => X"2326f100",
		16#23e7# => X"83270102",
		16#23e8# => X"93871700",
		16#23e9# => X"2320f102",
		16#23ea# => X"8327c100",
		16#23eb# => X"938707fe",
		16#23ec# => X"63f4fb00",
		16#23ed# => X"6f108028",
		16#23ee# => X"03270105",
		16#23ef# => X"93972700",
		16#23f0# => X"b387e700",
		16#23f1# => X"83a70700",
		16#23f2# => X"67800700",
		16#23f3# => X"13041400",
		16#23f4# => X"6ff01ff3",
		16#23f5# => X"b7470110",
		16#23f6# => X"93878791",
		16#23f7# => X"2322f104",
		16#23f8# => X"93770402",
		16#23f9# => X"63940700",
		16#23fa# => X"6f108008",
		16#23fb# => X"130c7c00",
		16#23fc# => X"137c8cff",
		16#23fd# => X"93078c00",
		16#23fe# => X"832c0c00",
		16#23ff# => X"032c4c00",
		16#2400# => X"232ef100",
		16#2401# => X"93771400",
		16#2402# => X"63800702",
		16#2403# => X"b3e78c01",
		16#2404# => X"638c0700",
		16#2405# => X"93070003",
		16#2406# => X"230cf10a",
		16#2407# => X"8347c100",
		16#2408# => X"13642400",
		16#2409# => X"a30cf10a",
		16#240a# => X"1374f4bf",
		16#240b# => X"93072000",
		16#240c# => X"6f00d06d",
		16#240d# => X"13050900",
		16#240e# => X"efd09f9f",
		16#240f# => X"83274500",
		16#2410# => X"13850700",
		16#2411# => X"232ef102",
		16#2412# => X"ef80cffc",
		16#2413# => X"232aa102",
		16#2414# => X"13050900",
		16#2415# => X"efd0df9d",
		16#2416# => X"83278500",
		16#2417# => X"232af100",
		16#2418# => X"83274103",
		16#2419# => X"e38407f2",
		16#241a# => X"83274101",
		16#241b# => X"e38007f2",
		16#241c# => X"83c70700",
		16#241d# => X"e38c07f0",
		16#241e# => X"13640440",
		16#241f# => X"6ff01ff1",
		16#2420# => X"8347710b",
		16#2421# => X"e39407f0",
		16#2422# => X"93070002",
		16#2423# => X"a30bf10a",
		16#2424# => X"6ff0dfef",
		16#2425# => X"13641400",
		16#2426# => X"6ff05fef",
		16#2427# => X"83270c00",
		16#2428# => X"130c4c00",
		16#2429# => X"2326f102",
		16#242a# => X"e3d207ee",
		16#242b# => X"b307f040",
		16#242c# => X"2326f102",
		16#242d# => X"13644400",
		16#242e# => X"6ff05fed",
		16#242f# => X"9307b002",
		16#2430# => X"6ff0dffc",
		16#2431# => X"83270102",
		16#2432# => X"1307a002",
		16#2433# => X"938c1700",
		16#2434# => X"83c70700",
		16#2435# => X"2326f100",
		16#2436# => X"6398e704",
		16#2437# => X"032b0c00",
		16#2438# => X"93074c00",
		16#2439# => X"63540b00",
		16#243a# => X"130bf0ff",
		16#243b# => X"138c0700",
		16#243c# => X"23209103",
		16#243d# => X"6ff09fe9",
		16#243e# => X"13050b00",
		16#243f# => X"9305a000",
		16#2440# => X"ef900053",
		16#2441# => X"938c1c00",
		16#2442# => X"83c7fcff",
		16#2443# => X"330bb501",
		16#2444# => X"2326f100",
		16#2445# => X"8327c100",
		16#2446# => X"938d07fd",
		16#2447# => X"e3febafd",
		16#2448# => X"23209103",
		16#2449# => X"6ff05fe8",
		16#244a# => X"130b0000",
		16#244b# => X"6ff09ffe",
		16#244c# => X"13640408",
		16#244d# => X"6ff09fe5",
		16#244e# => X"832c0102",
		16#244f# => X"23260102",
		16#2450# => X"0325c102",
		16#2451# => X"9305a000",
		16#2452# => X"938c1c00",
		16#2453# => X"ef90404e",
		16#2454# => X"8327c100",
		16#2455# => X"938707fd",
		16#2456# => X"b387a700",
		16#2457# => X"2326f102",
		16#2458# => X"83c7fcff",
		16#2459# => X"2326f100",
		16#245a# => X"938707fd",
		16#245b# => X"e3fafafc",
		16#245c# => X"6ff01ffb",
		16#245d# => X"13648400",
		16#245e# => X"6ff05fe1",
		16#245f# => X"83270102",
		16#2460# => X"03c70700",
		16#2461# => X"93078006",
		16#2462# => X"631cf700",
		16#2463# => X"83270102",
		16#2464# => X"13640420",
		16#2465# => X"93871700",
		16#2466# => X"2320f102",
		16#2467# => X"6ff01fdf",
		16#2468# => X"13640404",
		16#2469# => X"6ff09fde",
		16#246a# => X"83270102",
		16#246b# => X"03c70700",
		16#246c# => X"9307c006",
		16#246d# => X"631cf700",
		16#246e# => X"83270102",
		16#246f# => X"93871700",
		16#2470# => X"2320f102",
		16#2471# => X"13640402",
		16#2472# => X"6ff05fdc",
		16#2473# => X"13640401",
		16#2474# => X"6ff0dfdb",
		16#2475# => X"93074c00",
		16#2476# => X"232ef100",
		16#2477# => X"83270c00",
		16#2478# => X"a30b010a",
		16#2479# => X"230ef112",
		16#247a# => X"23280100",
		16#247b# => X"130b1000",
		16#247c# => X"930a0000",
		16#247d# => X"130c0000",
		16#247e# => X"930b0000",
		16#247f# => X"930c0000",
		16#2480# => X"9304c113",
		16#2481# => X"23285103",
		16#2482# => X"63d46a01",
		16#2483# => X"23286103",
		16#2484# => X"0347710b",
		16#2485# => X"63080700",
		16#2486# => X"83270103",
		16#2487# => X"93871700",
		16#2488# => X"2328f102",
		16#2489# => X"937d2400",
		16#248a# => X"63880d00",
		16#248b# => X"83270103",
		16#248c# => X"93872700",
		16#248d# => X"2328f102",
		16#248e# => X"93774408",
		16#248f# => X"2324f104",
		16#2490# => X"639c0706",
		16#2491# => X"8327c102",
		16#2492# => X"03270103",
		16#2493# => X"338ee740",
		16#2494# => X"6354c007",
		16#2495# => X"b74e0110",
		16#2496# => X"130f0001",
		16#2497# => X"938ece1c",
		16#2498# => X"930f7000",
		16#2499# => X"8326810d",
		16#249a# => X"2320dd01",
		16#249b# => X"0327c10d",
		16#249c# => X"93861600",
		16#249d# => X"13068d00",
		16#249e# => X"6354cf01",
		16#249f# => X"6f00d07d",
		16#24a0# => X"3307ee00",
		16#24a1# => X"2322cd01",
		16#24a2# => X"232ee10c",
		16#24a3# => X"232cd10c",
		16#24a4# => X"13077000",
		16#24a5# => X"130d0600",
		16#24a6# => X"6350d702",
		16#24a7# => X"1306410d",
		16#24a8# => X"93850900",
		16#24a9# => X"13050900",
		16#24aa# => X"ef209079",
		16#24ab# => X"63040500",
		16#24ac# => X"6f105022",
		16#24ad# => X"130dc10f",
		16#24ae# => X"0347710b",
		16#24af# => X"630a0704",
		16#24b0# => X"1307710b",
		16#24b1# => X"2320ed00",
		16#24b2# => X"13071000",
		16#24b3# => X"2322ed00",
		16#24b4# => X"0327c10d",
		16#24b5# => X"93067000",
		16#24b6# => X"130d8d00",
		16#24b7# => X"13071700",
		16#24b8# => X"232ee10c",
		16#24b9# => X"0327810d",
		16#24ba# => X"13071700",
		16#24bb# => X"232ce10c",
		16#24bc# => X"63d0e602",
		16#24bd# => X"1306410d",
		16#24be# => X"93850900",
		16#24bf# => X"13050900",
		16#24c0# => X"ef201074",
		16#24c1# => X"63040500",
		16#24c2# => X"6f10d01c",
		16#24c3# => X"130dc10f",
		16#24c4# => X"638a0d04",
		16#24c5# => X"1307810b",
		16#24c6# => X"2320ed00",
		16#24c7# => X"13072000",
		16#24c8# => X"2322ed00",
		16#24c9# => X"0327c10d",
		16#24ca# => X"93067000",
		16#24cb# => X"130d8d00",
		16#24cc# => X"13072700",
		16#24cd# => X"232ee10c",
		16#24ce# => X"0327810d",
		16#24cf# => X"13071700",
		16#24d0# => X"232ce10c",
		16#24d1# => X"63d0e602",
		16#24d2# => X"1306410d",
		16#24d3# => X"93850900",
		16#24d4# => X"13050900",
		16#24d5# => X"ef20d06e",
		16#24d6# => X"63040500",
		16#24d7# => X"6f109017",
		16#24d8# => X"130dc10f",
		16#24d9# => X"83278104",
		16#24da# => X"13070008",
		16#24db# => X"6398e706",
		16#24dc# => X"8327c102",
		16#24dd# => X"03270103",
		16#24de# => X"b38de740",
		16#24df# => X"6350b007",
		16#24e0# => X"93070001",
		16#24e1# => X"130e7000",
		16#24e2# => X"0327810d",
		16#24e3# => X"8326c10d",
		16#24e4# => X"13068d00",
		16#24e5# => X"13071700",
		16#24e6# => X"e3ccb771",
		16#24e7# => X"83278101",
		16#24e8# => X"2322bd01",
		16#24e9# => X"b38ddd00",
		16#24ea# => X"2320fd00",
		16#24eb# => X"232eb10d",
		16#24ec# => X"232ce10c",
		16#24ed# => X"93067000",
		16#24ee# => X"130d0600",
		16#24ef# => X"63d0e602",
		16#24f0# => X"1306410d",
		16#24f1# => X"93850900",
		16#24f2# => X"13050900",
		16#24f3# => X"ef205067",
		16#24f4# => X"63040500",
		16#24f5# => X"6f101010",
		16#24f6# => X"130dc10f",
		16#24f7# => X"b38a6a41",
		16#24f8# => X"63505007",
		16#24f9# => X"930d0001",
		16#24fa# => X"13087000",
		16#24fb# => X"83278101",
		16#24fc# => X"0327810d",
		16#24fd# => X"8326c10d",
		16#24fe# => X"2320fd00",
		16#24ff# => X"13071700",
		16#2500# => X"13068d00",
		16#2501# => X"e3ce5d6f",
		16#2502# => X"23225d01",
		16#2503# => X"b38ada00",
		16#2504# => X"232e510d",
		16#2505# => X"232ce10c",
		16#2506# => X"93067000",
		16#2507# => X"130d0600",
		16#2508# => X"63d0e602",
		16#2509# => X"1306410d",
		16#250a# => X"93850900",
		16#250b# => X"13050900",
		16#250c# => X"ef201061",
		16#250d# => X"63040500",
		16#250e# => X"6f10d009",
		16#250f# => X"130dc10f",
		16#2510# => X"13770410",
		16#2511# => X"832dc10d",
		16#2512# => X"e31c076e",
		16#2513# => X"8327810d",
		16#2514# => X"3303bb01",
		16#2515# => X"23209d00",
		16#2516# => X"93871700",
		16#2517# => X"23226d01",
		16#2518# => X"232e610c",
		16#2519# => X"232cf10c",
		16#251a# => X"13077000",
		16#251b# => X"130d8d00",
		16#251c# => X"6344f700",
		16#251d# => X"6f104019",
		16#251e# => X"1306410d",
		16#251f# => X"93850900",
		16#2520# => X"13050900",
		16#2521# => X"ef20d05b",
		16#2522# => X"63040500",
		16#2523# => X"6f109004",
		16#2524# => X"130dc10f",
		16#2525# => X"6f104017",
		16#2526# => X"13640401",
		16#2527# => X"93770402",
		16#2528# => X"638e0704",
		16#2529# => X"130c7c00",
		16#252a# => X"137c8cff",
		16#252b# => X"93078c00",
		16#252c# => X"832c0c00",
		16#252d# => X"032c4c00",
		16#252e# => X"232ef100",
		16#252f# => X"635e0c00",
		16#2530# => X"b30c9041",
		16#2531# => X"b3379001",
		16#2532# => X"330c8041",
		16#2533# => X"330cfc40",
		16#2534# => X"9307d002",
		16#2535# => X"a30bf10a",
		16#2536# => X"9307f0ff",
		16#2537# => X"e318fb3c",
		16#2538# => X"e31a0c44",
		16#2539# => X"93079000",
		16#253a# => X"e3e69745",
		16#253b# => X"938c0c03",
		16#253c# => X"a30f9119",
		16#253d# => X"9304f119",
		16#253e# => X"6f005041",
		16#253f# => X"93074c00",
		16#2540# => X"232ef100",
		16#2541# => X"93770401",
		16#2542# => X"63880700",
		16#2543# => X"832c0c00",
		16#2544# => X"13dcfc41",
		16#2545# => X"6ff09ffa",
		16#2546# => X"93770404",
		16#2547# => X"832c0c00",
		16#2548# => X"63880700",
		16#2549# => X"939c0c01",
		16#254a# => X"93dc0c41",
		16#254b# => X"6ff05ffe",
		16#254c# => X"93770420",
		16#254d# => X"e38e07fc",
		16#254e# => X"939c8c01",
		16#254f# => X"93dc8c41",
		16#2550# => X"6ff01ffd",
		16#2551# => X"93778400",
		16#2552# => X"638a070a",
		16#2553# => X"93074c00",
		16#2554# => X"232ef100",
		16#2555# => X"83270c00",
		16#2556# => X"03a60700",
		16#2557# => X"83a64700",
		16#2558# => X"03a78700",
		16#2559# => X"83a7c700",
		16#255a# => X"2320c10e",
		16#255b# => X"2322d10e",
		16#255c# => X"2324e10e",
		16#255d# => X"1305010e",
		16#255e# => X"2326f10e",
		16#255f# => X"efd08fc4",
		16#2560# => X"232ea10a",
		16#2561# => X"93072000",
		16#2562# => X"6310f50c",
		16#2563# => X"8327010e",
		16#2564# => X"93050109",
		16#2565# => X"1305010a",
		16#2566# => X"2320f10a",
		16#2567# => X"8327410e",
		16#2568# => X"23280108",
		16#2569# => X"232a0108",
		16#256a# => X"2322f10a",
		16#256b# => X"8327810e",
		16#256c# => X"232c0108",
		16#256d# => X"232e0108",
		16#256e# => X"2324f10a",
		16#256f# => X"8327c10e",
		16#2570# => X"2326f10a",
		16#2571# => X"ef501052",
		16#2572# => X"63560500",
		16#2573# => X"9307d002",
		16#2574# => X"a30bf10a",
		16#2575# => X"0327c100",
		16#2576# => X"93077004",
		16#2577# => X"63c0e706",
		16#2578# => X"b7440110",
		16#2579# => X"9384448f",
		16#257a# => X"1374f4f7",
		16#257b# => X"23280100",
		16#257c# => X"130b3000",
		16#257d# => X"930a0000",
		16#257e# => X"6f005032",
		16#257f# => X"130c7c00",
		16#2580# => X"137c8cff",
		16#2581# => X"83250c00",
		16#2582# => X"03264c00",
		16#2583# => X"93078c00",
		16#2584# => X"1305010a",
		16#2585# => X"232ef100",
		16#2586# => X"ef801027",
		16#2587# => X"8327010a",
		16#2588# => X"2320f10e",
		16#2589# => X"8327410a",
		16#258a# => X"2322f10e",
		16#258b# => X"8327810a",
		16#258c# => X"2324f10e",
		16#258d# => X"8327c10a",
		16#258e# => X"6ff0dff3",
		16#258f# => X"b7440110",
		16#2590# => X"9384848f",
		16#2591# => X"6ff05ffa",
		16#2592# => X"93071000",
		16#2593# => X"631cf502",
		16#2594# => X"8327c10e",
		16#2595# => X"63d60700",
		16#2596# => X"9307d002",
		16#2597# => X"a30bf10a",
		16#2598# => X"0327c100",
		16#2599# => X"93077004",
		16#259a# => X"63c8e700",
		16#259b# => X"b7440110",
		16#259c# => X"9384c48f",
		16#259d# => X"6ff05ff7",
		16#259e# => X"b7440110",
		16#259f# => X"93840490",
		16#25a0# => X"6ff09ff6",
		16#25a1# => X"8327c100",
		16#25a2# => X"93fbf7fd",
		16#25a3# => X"93071004",
		16#25a4# => X"639efb08",
		16#25a5# => X"8326c100",
		16#25a6# => X"93070003",
		16#25a7# => X"230cf10a",
		16#25a8# => X"13071006",
		16#25a9# => X"93078005",
		16#25aa# => X"6394e600",
		16#25ab# => X"93078007",
		16#25ac# => X"a30cf10a",
		16#25ad# => X"93073006",
		16#25ae# => X"13642400",
		16#25af# => X"63dc674d",
		16#25b0# => X"93051b00",
		16#25b1# => X"13050900",
		16#25b2# => X"efd00fdf",
		16#25b3# => X"93040500",
		16#25b4# => X"6318054c",
		16#25b5# => X"83d7c900",
		16#25b6# => X"93e70704",
		16#25b7# => X"2396f900",
		16#25b8# => X"83d7c900",
		16#25b9# => X"93f70704",
		16#25ba# => X"639a07fa",
		16#25bb# => X"8320c11d",
		16#25bc# => X"0324811d",
		16#25bd# => X"03258102",
		16#25be# => X"8324411d",
		16#25bf# => X"0329011d",
		16#25c0# => X"8329c11c",
		16#25c1# => X"032a811c",
		16#25c2# => X"832a411c",
		16#25c3# => X"032b011c",
		16#25c4# => X"832bc11b",
		16#25c5# => X"032c811b",
		16#25c6# => X"832c411b",
		16#25c7# => X"032d011b",
		16#25c8# => X"832dc11a",
		16#25c9# => X"1301011e",
		16#25ca# => X"67800000",
		16#25cb# => X"9307f0ff",
		16#25cc# => X"630cfb46",
		16#25cd# => X"93077004",
		16#25ce# => X"23280100",
		16#25cf# => X"6394fb00",
		16#25d0# => X"630a0b46",
		16#25d1# => X"832ac10e",
		16#25d2# => X"93670410",
		16#25d3# => X"2328f102",
		16#25d4# => X"23240104",
		16#25d5# => X"032e010e",
		16#25d6# => X"832d410e",
		16#25d7# => X"832c810e",
		16#25d8# => X"63da0a00",
		16#25d9# => X"b7070080",
		16#25da# => X"b3ca5701",
		16#25db# => X"9307d002",
		16#25dc# => X"2324f104",
		16#25dd# => X"93071004",
		16#25de# => X"6398fb48",
		16#25df# => X"1305010a",
		16#25e0# => X"2320c10b",
		16#25e1# => X"2324910b",
		16#25e2# => X"2322b10b",
		16#25e3# => X"2326510b",
		16#25e4# => X"ef809034",
		16#25e5# => X"1306c10b",
		16#25e6# => X"eff0cfb3",
		16#25e7# => X"13860500",
		16#25e8# => X"93050500",
		16#25e9# => X"1305010a",
		16#25ea# => X"ef80100e",
		16#25eb# => X"8327010a",
		16#25ec# => X"13060107",
		16#25ed# => X"93050108",
		16#25ee# => X"2320f108",
		16#25ef# => X"8327410a",
		16#25f0# => X"13050109",
		16#25f1# => X"23280106",
		16#25f2# => X"2322f108",
		16#25f3# => X"8327810a",
		16#25f4# => X"232a0106",
		16#25f5# => X"232c0106",
		16#25f6# => X"2324f108",
		16#25f7# => X"8327c10a",
		16#25f8# => X"2326f108",
		16#25f9# => X"b707fc3f",
		16#25fa# => X"232ef106",
		16#25fb# => X"ef509045",
		16#25fc# => X"03280109",
		16#25fd# => X"03264109",
		16#25fe# => X"83268109",
		16#25ff# => X"832cc109",
		16#2600# => X"93050109",
		16#2601# => X"1305010a",
		16#2602# => X"2320010b",
		16#2603# => X"232c0105",
		16#2604# => X"2322c10a",
		16#2605# => X"232ac104",
		16#2606# => X"2324d10a",
		16#2607# => X"2326d104",
		16#2608# => X"2326910b",
		16#2609# => X"23280108",
		16#260a# => X"232a0108",
		16#260b# => X"232c0108",
		16#260c# => X"232e0108",
		16#260d# => X"ef505008",
		16#260e# => X"8326c104",
		16#260f# => X"03264105",
		16#2610# => X"03288105",
		16#2611# => X"63160500",
		16#2612# => X"13071000",
		16#2613# => X"232ee10a",
		16#2614# => X"8327c100",
		16#2615# => X"13071006",
		16#2616# => X"6394e736",
		16#2617# => X"374a0110",
		16#2618# => X"130a4a90",
		16#2619# => X"130efbff",
		16#261a# => X"938d0400",
		16#261b# => X"b7070340",
		16#261c# => X"93050109",
		16#261d# => X"232ac108",
		16#261e# => X"1305010a",
		16#261f# => X"13060108",
		16#2620# => X"232cc105",
		16#2621# => X"23280109",
		16#2622# => X"2326f108",
		16#2623# => X"232cd108",
		16#2624# => X"232e9109",
		16#2625# => X"23200108",
		16#2626# => X"23220108",
		16#2627# => X"23240108",
		16#2628# => X"ef50503a",
		16#2629# => X"0326010a",
		16#262a# => X"8326410a",
		16#262b# => X"1305010a",
		16#262c# => X"232ac104",
		16#262d# => X"2326d104",
		16#262e# => X"ef80c04e",
		16#262f# => X"93050500",
		16#2630# => X"930a0500",
		16#2631# => X"1305010a",
		16#2632# => X"832c810a",
		16#2633# => X"032cc10a",
		16#2634# => X"ef808063",
		16#2635# => X"8327010a",
		16#2636# => X"03264105",
		16#2637# => X"8326c104",
		16#2638# => X"2328f106",
		16#2639# => X"8327410a",
		16#263a# => X"2320c108",
		16#263b# => X"93050108",
		16#263c# => X"232af106",
		16#263d# => X"8327810a",
		16#263e# => X"13060107",
		16#263f# => X"13050109",
		16#2640# => X"232cf106",
		16#2641# => X"8327c10a",
		16#2642# => X"23249109",
		16#2643# => X"23268109",
		16#2644# => X"232ef106",
		16#2645# => X"2322d108",
		16#2646# => X"ef609078",
		16#2647# => X"b3055a01",
		16#2648# => X"83c50500",
		16#2649# => X"032e8105",
		16#264a# => X"032cc109",
		16#264b# => X"938d1d00",
		16#264c# => X"83220109",
		16#264d# => X"832f4109",
		16#264e# => X"032f8109",
		16#264f# => X"2326c105",
		16#2650# => X"a38fbdfe",
		16#2651# => X"9307f0ff",
		16#2652# => X"930c0c00",
		16#2653# => X"6308fe06",
		16#2654# => X"130efeff",
		16#2655# => X"93050109",
		16#2656# => X"1305010a",
		16#2657# => X"2326e107",
		16#2658# => X"2324f107",
		16#2659# => X"23225106",
		16#265a# => X"2320c107",
		16#265b# => X"2320510a",
		16#265c# => X"232e5104",
		16#265d# => X"2322f10b",
		16#265e# => X"232cf105",
		16#265f# => X"2324e10b",
		16#2660# => X"232ae105",
		16#2661# => X"2326810b",
		16#2662# => X"23280108",
		16#2663# => X"232a0108",
		16#2664# => X"232c0108",
		16#2665# => X"232e0108",
		16#2666# => X"ef500072",
		16#2667# => X"83264105",
		16#2668# => X"03268105",
		16#2669# => X"0328c105",
		16#266a# => X"032e0106",
		16#266b# => X"83224106",
		16#266c# => X"832f8106",
		16#266d# => X"032fc106",
		16#266e# => X"e31a05ea",
		16#266f# => X"b70cfe3f",
		16#2670# => X"93050109",
		16#2671# => X"1305010a",
		16#2672# => X"2320510a",
		16#2673# => X"232e5104",
		16#2674# => X"2322f10b",
		16#2675# => X"232cf105",
		16#2676# => X"2324e10b",
		16#2677# => X"232ae105",
		16#2678# => X"2326810b",
		16#2679# => X"23280108",
		16#267a# => X"232a0108",
		16#267b# => X"232c0108",
		16#267c# => X"232e9109",
		16#267d# => X"ef500079",
		16#267e# => X"6344a004",
		16#267f# => X"8322c105",
		16#2680# => X"832f8105",
		16#2681# => X"032f4105",
		16#2682# => X"93050109",
		16#2683# => X"1305010a",
		16#2684# => X"2320510a",
		16#2685# => X"2322f10b",
		16#2686# => X"2324e10b",
		16#2687# => X"2326810b",
		16#2688# => X"23280108",
		16#2689# => X"232a0108",
		16#268a# => X"232c0108",
		16#268b# => X"232e9109",
		16#268c# => X"ef508068",
		16#268d# => X"6310051c",
		16#268e# => X"93fa1a00",
		16#268f# => X"638c0a1a",
		16#2690# => X"0346fa00",
		16#2691# => X"2326b10d",
		16#2692# => X"93050003",
		16#2693# => X"8326c10c",
		16#2694# => X"9387f6ff",
		16#2695# => X"2326f10c",
		16#2696# => X"83c7f6ff",
		16#2697# => X"6388c716",
		16#2698# => X"13069003",
		16#2699# => X"6398c716",
		16#269a# => X"8347aa00",
		16#269b# => X"a38ff6fe",
		16#269c# => X"138a0d00",
		16#269d# => X"13077004",
		16#269e# => X"330a9a40",
		16#269f# => X"832cc10b",
		16#26a0# => X"639aeb2a",
		16#26a1# => X"1307d0ff",
		16#26a2# => X"63c4ec00",
		16#26a3# => X"63589b33",
		16#26a4# => X"8327c100",
		16#26a5# => X"9387e7ff",
		16#26a6# => X"2326f100",
		16#26a7# => X"8327c100",
		16#26a8# => X"938afcff",
		16#26a9# => X"232e510b",
		16#26aa# => X"93f6f7fd",
		16#26ab# => X"93051004",
		16#26ac# => X"0347c100",
		16#26ad# => X"13060000",
		16#26ae# => X"6398b600",
		16#26af# => X"1307f700",
		16#26b0# => X"1377f70f",
		16#26b1# => X"13061000",
		16#26b2# => X"2302e10c",
		16#26b3# => X"9307b002",
		16#26b4# => X"63d80a00",
		16#26b5# => X"930a1000",
		16#26b6# => X"b38a9a41",
		16#26b7# => X"9307d002",
		16#26b8# => X"a302f10c",
		16#26b9# => X"93079000",
		16#26ba# => X"63dc5729",
		16#26bb# => X"930b310d",
		16#26bc# => X"938c0b00",
		16#26bd# => X"930d9000",
		16#26be# => X"9305a000",
		16#26bf# => X"13850a00",
		16#26c0# => X"ef80903d",
		16#26c1# => X"13050503",
		16#26c2# => X"a38fabfe",
		16#26c3# => X"9305a000",
		16#26c4# => X"13850a00",
		16#26c5# => X"ef801034",
		16#26c6# => X"138cfbff",
		16#26c7# => X"930a0500",
		16#26c8# => X"63c2ad24",
		16#26c9# => X"930a0503",
		16#26ca# => X"938bebff",
		16#26cb# => X"a30f5cff",
		16#26cc# => X"9307610c",
		16#26cd# => X"63ec9b23",
		16#26ce# => X"1307410c",
		16#26cf# => X"b387e740",
		16#26d0# => X"2320f104",
		16#26d1# => X"338b4701",
		16#26d2# => X"93071000",
		16#26d3# => X"63c64701",
		16#26d4# => X"93771400",
		16#26d5# => X"63860700",
		16#26d6# => X"83274102",
		16#26d7# => X"330bfb00",
		16#26d8# => X"1374f4bf",
		16#26d9# => X"93670410",
		16#26da# => X"2328f102",
		16#26db# => X"130c0000",
		16#26dc# => X"930b0000",
		16#26dd# => X"930c0000",
		16#26de# => X"83278104",
		16#26df# => X"63860700",
		16#26e0# => X"1307d002",
		16#26e1# => X"a30be10a",
		16#26e2# => X"03240103",
		16#26e3# => X"930a0000",
		16#26e4# => X"6ff04fe7",
		16#26e5# => X"23280100",
		16#26e6# => X"9304c113",
		16#26e7# => X"6ff09fba",
		16#26e8# => X"2328a100",
		16#26e9# => X"6ff01fba",
		16#26ea# => X"23280100",
		16#26eb# => X"130b6000",
		16#26ec# => X"6ff05fb9",
		16#26ed# => X"23286101",
		16#26ee# => X"130b1000",
		16#26ef# => X"6ff09fb8",
		16#26f0# => X"374a0110",
		16#26f1# => X"130a8a91",
		16#26f2# => X"6ff0dfc9",
		16#26f3# => X"a38fb6fe",
		16#26f4# => X"6ff0dfe7",
		16#26f5# => X"93871700",
		16#26f6# => X"93f7f70f",
		16#26f7# => X"6ff01fe9",
		16#26f8# => X"130a1a00",
		16#26f9# => X"a30feafe",
		16#26fa# => X"b3074c41",
		16#26fb# => X"e3da07fe",
		16#26fc# => X"6ff05fe8",
		16#26fd# => X"8327c104",
		16#26fe# => X"138a0d00",
		16#26ff# => X"13070003",
		16#2700# => X"338cfd00",
		16#2701# => X"6ff05ffe",
		16#2702# => X"93076004",
		16#2703# => X"638efb00",
		16#2704# => X"93075004",
		16#2705# => X"130c1b00",
		16#2706# => X"6384fb00",
		16#2707# => X"130c0b00",
		16#2708# => X"13062000",
		16#2709# => X"6f00c000",
		16#270a# => X"130c0b00",
		16#270b# => X"13063000",
		16#270c# => X"9307010c",
		16#270d# => X"1308c10c",
		16#270e# => X"1307c10b",
		16#270f# => X"93060c00",
		16#2710# => X"9305010a",
		16#2711# => X"13050900",
		16#2712# => X"2320c10b",
		16#2713# => X"2326c105",
		16#2714# => X"2322b10b",
		16#2715# => X"2324910b",
		16#2716# => X"2326510b",
		16#2717# => X"efc04f91",
		16#2718# => X"93077004",
		16#2719# => X"93040500",
		16#271a# => X"032ec104",
		16#271b# => X"6396fb00",
		16#271c# => X"93771400",
		16#271d# => X"6380070a",
		16#271e# => X"93076004",
		16#271f# => X"338a8401",
		16#2720# => X"639efb04",
		16#2721# => X"03c70400",
		16#2722# => X"93070003",
		16#2723# => X"6314f704",
		16#2724# => X"93050109",
		16#2725# => X"1305010a",
		16#2726# => X"2320c10b",
		16#2727# => X"2326c105",
		16#2728# => X"2322b10b",
		16#2729# => X"2324910b",
		16#272a# => X"2326510b",
		16#272b# => X"23280108",
		16#272c# => X"232a0108",
		16#272d# => X"232c0108",
		16#272e# => X"232e0108",
		16#272f# => X"ef50c03f",
		16#2730# => X"032ec104",
		16#2731# => X"63080500",
		16#2732# => X"93071000",
		16#2733# => X"338c8741",
		16#2734# => X"232e810b",
		16#2735# => X"8327c10b",
		16#2736# => X"330afa00",
		16#2737# => X"93050109",
		16#2738# => X"1305010a",
		16#2739# => X"2320c10b",
		16#273a# => X"2322b10b",
		16#273b# => X"2324910b",
		16#273c# => X"2326510b",
		16#273d# => X"23280108",
		16#273e# => X"232a0108",
		16#273f# => X"232c0108",
		16#2740# => X"232e0108",
		16#2741# => X"ef50403b",
		16#2742# => X"13070003",
		16#2743# => X"631e0500",
		16#2744# => X"2326410d",
		16#2745# => X"032ac10c",
		16#2746# => X"6ff0dfd5",
		16#2747# => X"93861700",
		16#2748# => X"2326d10c",
		16#2749# => X"2380e700",
		16#274a# => X"8327c10c",
		16#274b# => X"e3e847ff",
		16#274c# => X"6ff05ffe",
		16#274d# => X"13076004",
		16#274e# => X"e392ebd6",
		16#274f# => X"63549007",
		16#2750# => X"63160b00",
		16#2751# => X"13771400",
		16#2752# => X"6306070c",
		16#2753# => X"83274102",
		16#2754# => X"3387fc00",
		16#2755# => X"330beb00",
		16#2756# => X"93076006",
		16#2757# => X"2326f100",
		16#2758# => X"6f008009",
		16#2759# => X"930b0c00",
		16#275a# => X"6ff01fd9",
		16#275b# => X"938b1b00",
		16#275c# => X"03c7fbff",
		16#275d# => X"93871700",
		16#275e# => X"a38fe7fe",
		16#275f# => X"6ff09fdb",
		16#2760# => X"1307610c",
		16#2761# => X"63180600",
		16#2762# => X"93070003",
		16#2763# => X"2303f10c",
		16#2764# => X"1307710c",
		16#2765# => X"938a0a03",
		16#2766# => X"93071700",
		16#2767# => X"23005701",
		16#2768# => X"6ff09fd9",
		16#2769# => X"63160b00",
		16#276a# => X"13771400",
		16#276b# => X"63080706",
		16#276c# => X"83274102",
		16#276d# => X"13871700",
		16#276e# => X"6ff0dff9",
		16#276f# => X"63c04c03",
		16#2770# => X"13771400",
		16#2771# => X"138b0c00",
		16#2772# => X"63060700",
		16#2773# => X"83274102",
		16#2774# => X"338bfc00",
		16#2775# => X"93077006",
		16#2776# => X"6ff05ff8",
		16#2777# => X"83274102",
		16#2778# => X"330bfa00",
		16#2779# => X"93077006",
		16#277a# => X"2326f100",
		16#277b# => X"63469001",
		16#277c# => X"33039b41",
		16#277d# => X"130b1300",
		16#277e# => X"937b0440",
		16#277f# => X"130c0000",
		16#2780# => X"e38c0bd6",
		16#2781# => X"930b0000",
		16#2782# => X"e35890d7",
		16#2783# => X"9306f00f",
		16#2784# => X"6f00c003",
		16#2785# => X"138b0c00",
		16#2786# => X"6ff01ff4",
		16#2787# => X"93076006",
		16#2788# => X"2326f100",
		16#2789# => X"130b1000",
		16#278a# => X"6ff01ffd",
		16#278b# => X"63569703",
		16#278c# => X"83274101",
		16#278d# => X"b38cec40",
		16#278e# => X"03c71700",
		16#278f# => X"63080702",
		16#2790# => X"93871700",
		16#2791# => X"938b1b00",
		16#2792# => X"232af100",
		16#2793# => X"83274101",
		16#2794# => X"03c70700",
		16#2795# => X"e31cd7fc",
		16#2796# => X"83254103",
		16#2797# => X"33858b01",
		16#2798# => X"ef80007d",
		16#2799# => X"330b6501",
		16#279a# => X"6ff01fd1",
		16#279b# => X"130c1c00",
		16#279c# => X"6ff0dffd",
		16#279d# => X"13074c00",
		16#279e# => X"232ee100",
		16#279f# => X"13770402",
		16#27a0# => X"83270c00",
		16#27a1# => X"63000702",
		16#27a2# => X"03278102",
		16#27a3# => X"23a0e700",
		16#27a4# => X"1357f741",
		16#27a5# => X"23a2e700",
		16#27a6# => X"032cc101",
		16#27a7# => X"83240102",
		16#27a8# => X"6ff08f85",
		16#27a9# => X"13770401",
		16#27aa# => X"63080700",
		16#27ab# => X"03278102",
		16#27ac# => X"23a0e700",
		16#27ad# => X"6ff05ffe",
		16#27ae# => X"13770404",
		16#27af# => X"63080700",
		16#27b0# => X"03578102",
		16#27b1# => X"2390e700",
		16#27b2# => X"6ff01ffd",
		16#27b3# => X"13740420",
		16#27b4# => X"e30e04fc",
		16#27b5# => X"03478102",
		16#27b6# => X"2380e700",
		16#27b7# => X"6ff0dffb",
		16#27b8# => X"13640401",
		16#27b9# => X"93770402",
		16#27ba# => X"63880704",
		16#27bb# => X"130c7c00",
		16#27bc# => X"137c8cff",
		16#27bd# => X"93078c00",
		16#27be# => X"832c0c00",
		16#27bf# => X"032c4c00",
		16#27c0# => X"232ef100",
		16#27c1# => X"1374f4bf",
		16#27c2# => X"93070000",
		16#27c3# => X"a30b010a",
		16#27c4# => X"1307f0ff",
		16#27c5# => X"6302eb1a",
		16#27c6# => X"13070400",
		16#27c7# => X"b3e68c01",
		16#27c8# => X"1374f4f7",
		16#27c9# => X"639a0618",
		16#27ca# => X"630c0b2e",
		16#27cb# => X"13071000",
		16#27cc# => X"6398e718",
		16#27cd# => X"6ff08fdb",
		16#27ce# => X"93074c00",
		16#27cf# => X"232ef100",
		16#27d0# => X"93770401",
		16#27d1# => X"63860700",
		16#27d2# => X"832c0c00",
		16#27d3# => X"6f000001",
		16#27d4# => X"93770404",
		16#27d5# => X"63880700",
		16#27d6# => X"835c0c00",
		16#27d7# => X"130c0000",
		16#27d8# => X"6ff05ffa",
		16#27d9# => X"93770420",
		16#27da# => X"e38007fe",
		16#27db# => X"834c0c00",
		16#27dc# => X"6ff0dffe",
		16#27dd# => X"93074c00",
		16#27de# => X"232ef100",
		16#27df# => X"b787ffff",
		16#27e0# => X"93c70783",
		16#27e1# => X"231cf10a",
		16#27e2# => X"b7470110",
		16#27e3# => X"93874790",
		16#27e4# => X"13078007",
		16#27e5# => X"832c0c00",
		16#27e6# => X"2322f104",
		16#27e7# => X"130c0000",
		16#27e8# => X"13642400",
		16#27e9# => X"93072000",
		16#27ea# => X"2326e100",
		16#27eb# => X"6ff01ff6",
		16#27ec# => X"93074c00",
		16#27ed# => X"232ef100",
		16#27ee# => X"a30b010a",
		16#27ef# => X"9307f0ff",
		16#27f0# => X"83240c00",
		16#27f1# => X"6304fb02",
		16#27f2# => X"13060b00",
		16#27f3# => X"93050000",
		16#27f4# => X"13850400",
		16#27f5# => X"efd08fba",
		16#27f6# => X"2328a100",
		16#27f7# => X"630c05e0",
		16#27f8# => X"330b9540",
		16#27f9# => X"23280100",
		16#27fa# => X"6ff0cfe0",
		16#27fb# => X"13850400",
		16#27fc# => X"ef705f82",
		16#27fd# => X"130b0500",
		16#27fe# => X"6ff0dffe",
		16#27ff# => X"13640401",
		16#2800# => X"93770402",
		16#2801# => X"63820702",
		16#2802# => X"130c7c00",
		16#2803# => X"137c8cff",
		16#2804# => X"93078c00",
		16#2805# => X"832c0c00",
		16#2806# => X"032c4c00",
		16#2807# => X"232ef100",
		16#2808# => X"93071000",
		16#2809# => X"6ff09fee",
		16#280a# => X"93074c00",
		16#280b# => X"232ef100",
		16#280c# => X"93770401",
		16#280d# => X"63860700",
		16#280e# => X"832c0c00",
		16#280f# => X"6f000001",
		16#2810# => X"93770404",
		16#2811# => X"63880700",
		16#2812# => X"835c0c00",
		16#2813# => X"130c0000",
		16#2814# => X"6ff01ffd",
		16#2815# => X"93770420",
		16#2816# => X"e38007fe",
		16#2817# => X"834c0c00",
		16#2818# => X"6ff0dffe",
		16#2819# => X"b7470110",
		16#281a# => X"93874790",
		16#281b# => X"6fe01ff7",
		16#281c# => X"93074c00",
		16#281d# => X"232ef100",
		16#281e# => X"93770401",
		16#281f# => X"63860700",
		16#2820# => X"832c0c00",
		16#2821# => X"6f000001",
		16#2822# => X"93770404",
		16#2823# => X"63880700",
		16#2824# => X"835c0c00",
		16#2825# => X"130c0000",
		16#2826# => X"6fe0dff6",
		16#2827# => X"93770420",
		16#2828# => X"e38007fe",
		16#2829# => X"834c0c00",
		16#282a# => X"6ff0dffe",
		16#282b# => X"13070400",
		16#282c# => X"93071000",
		16#282d# => X"6ff09fe6",
		16#282e# => X"13071000",
		16#282f# => X"6382e7c2",
		16#2830# => X"13072000",
		16#2831# => X"6382e712",
		16#2832# => X"9307011a",
		16#2833# => X"9316dc01",
		16#2834# => X"13f77c00",
		16#2835# => X"93dc3c00",
		16#2836# => X"13070703",
		16#2837# => X"b3ec9601",
		16#2838# => X"135c3c00",
		16#2839# => X"a38fe7fe",
		16#283a# => X"b3e68c01",
		16#283b# => X"9384f7ff",
		16#283c# => X"639e0602",
		16#283d# => X"93761400",
		16#283e# => X"638a0600",
		16#283f# => X"93060003",
		16#2840# => X"6306d700",
		16#2841# => X"a38fd4fe",
		16#2842# => X"9384e7ff",
		16#2843# => X"9307011a",
		16#2844# => X"930a0b00",
		16#2845# => X"23280100",
		16#2846# => X"338b9740",
		16#2847# => X"130c0000",
		16#2848# => X"930b0000",
		16#2849# => X"930c0000",
		16#284a# => X"6ff0cf8d",
		16#284b# => X"93870400",
		16#284c# => X"6ff0dff9",
		16#284d# => X"130a0000",
		16#284e# => X"930d011a",
		16#284f# => X"937a0440",
		16#2850# => X"930b9000",
		16#2851# => X"1306a000",
		16#2852# => X"93060000",
		16#2853# => X"13850c00",
		16#2854# => X"93050c00",
		16#2855# => X"ef30d036",
		16#2856# => X"13050503",
		16#2857# => X"a38fadfe",
		16#2858# => X"9384fdff",
		16#2859# => X"130a1a00",
		16#285a# => X"638a0a04",
		16#285b# => X"83274101",
		16#285c# => X"83c70700",
		16#285d# => X"6314fa04",
		16#285e# => X"9307f00f",
		16#285f# => X"6300fa04",
		16#2860# => X"63140c00",
		16#2861# => X"63fc9b03",
		16#2862# => X"83274103",
		16#2863# => X"8325c103",
		16#2864# => X"130a0000",
		16#2865# => X"b384f440",
		16#2866# => X"13860700",
		16#2867# => X"13850400",
		16#2868# => X"efe01fc1",
		16#2869# => X"83274101",
		16#286a# => X"83c71700",
		16#286b# => X"63880700",
		16#286c# => X"83274101",
		16#286d# => X"93871700",
		16#286e# => X"232af100",
		16#286f# => X"13850c00",
		16#2870# => X"93050c00",
		16#2871# => X"1306a000",
		16#2872# => X"93060000",
		16#2873# => X"ef308051",
		16#2874# => X"138c0500",
		16#2875# => X"b3e5a500",
		16#2876# => X"930c0500",
		16#2877# => X"e38805f2",
		16#2878# => X"938d0400",
		16#2879# => X"6ff01ff6",
		16#287a# => X"9304011a",
		16#287b# => X"03274104",
		16#287c# => X"93f7fc00",
		16#287d# => X"9384f4ff",
		16#287e# => X"b307f700",
		16#287f# => X"83c70700",
		16#2880# => X"93dc4c00",
		16#2881# => X"2380f400",
		16#2882# => X"9317cc01",
		16#2883# => X"b3ec9701",
		16#2884# => X"135c4c00",
		16#2885# => X"b3e78c01",
		16#2886# => X"e39a07fc",
		16#2887# => X"6ff01fef",
		16#2888# => X"9304011a",
		16#2889# => X"e39407ee",
		16#288a# => X"13771700",
		16#288b# => X"e30007ee",
		16#288c# => X"93070003",
		16#288d# => X"a30ff118",
		16#288e# => X"6ff0cfab",
		16#288f# => X"8327c100",
		16#2890# => X"e38c072e",
		16#2891# => X"8347c100",
		16#2892# => X"a30b010a",
		16#2893# => X"232e8101",
		16#2894# => X"230ef112",
		16#2895# => X"6fe05ff9",
		16#2896# => X"13070701",
		16#2897# => X"2322ed01",
		16#2898# => X"232ee10c",
		16#2899# => X"232cd10c",
		16#289a# => X"63dedf02",
		16#289b# => X"1306410d",
		16#289c# => X"93850900",
		16#289d# => X"13050900",
		16#289e# => X"232ef105",
		16#289f# => X"232cd105",
		16#28a0# => X"232ae105",
		16#28a1# => X"2326c105",
		16#28a2# => X"ef10907b",
		16#28a3# => X"e3140524",
		16#28a4# => X"832fc105",
		16#28a5# => X"832e8105",
		16#28a6# => X"032f4105",
		16#28a7# => X"032ec104",
		16#28a8# => X"1306c10f",
		16#28a9# => X"130e0eff",
		16#28aa# => X"130d0600",
		16#28ab# => X"6fe09ffb",
		16#28ac# => X"83258101",
		16#28ad# => X"93860601",
		16#28ae# => X"2322fd00",
		16#28af# => X"2320bd00",
		16#28b0# => X"232ed10c",
		16#28b1# => X"232ce10c",
		16#28b2# => X"6356ee02",
		16#28b3# => X"1306410d",
		16#28b4# => X"93850900",
		16#28b5# => X"13050900",
		16#28b6# => X"2326c105",
		16#28b7# => X"2324f104",
		16#28b8# => X"ef101076",
		16#28b9# => X"e318051e",
		16#28ba# => X"032ec104",
		16#28bb# => X"83278104",
		16#28bc# => X"1306c10f",
		16#28bd# => X"938d0dff",
		16#28be# => X"130d0600",
		16#28bf# => X"6ff0cf88",
		16#28c0# => X"93860601",
		16#28c1# => X"2322bd01",
		16#28c2# => X"232ed10c",
		16#28c3# => X"232ce10c",
		16#28c4# => X"6352e802",
		16#28c5# => X"1306410d",
		16#28c6# => X"93850900",
		16#28c7# => X"13050900",
		16#28c8# => X"23240105",
		16#28c9# => X"ef10d071",
		16#28ca# => X"e316051a",
		16#28cb# => X"03288104",
		16#28cc# => X"1306c10f",
		16#28cd# => X"938a0aff",
		16#28ce# => X"130d0600",
		16#28cf# => X"6ff00f8b",
		16#28d0# => X"8327c100",
		16#28d1# => X"13075006",
		16#28d2# => X"6354f772",
		16#28d3# => X"0327010e",
		16#28d4# => X"93050109",
		16#28d5# => X"1305010a",
		16#28d6# => X"2320e10a",
		16#28d7# => X"0327410e",
		16#28d8# => X"23280108",
		16#28d9# => X"232a0108",
		16#28da# => X"2322e10a",
		16#28db# => X"0327810e",
		16#28dc# => X"232c0108",
		16#28dd# => X"232e0108",
		16#28de# => X"2324e10a",
		16#28df# => X"0327c10e",
		16#28e0# => X"2326e10a",
		16#28e1# => X"ef405053",
		16#28e2# => X"631a0512",
		16#28e3# => X"b7470110",
		16#28e4# => X"9387c792",
		16#28e5# => X"2320fd00",
		16#28e6# => X"93071000",
		16#28e7# => X"2322fd00",
		16#28e8# => X"8327810d",
		16#28e9# => X"938d1d00",
		16#28ea# => X"232eb10d",
		16#28eb# => X"93871700",
		16#28ec# => X"232cf10c",
		16#28ed# => X"13077000",
		16#28ee# => X"130d8d00",
		16#28ef# => X"635ef700",
		16#28f0# => X"1306410d",
		16#28f1# => X"93850900",
		16#28f2# => X"13050900",
		16#28f3# => X"ef105067",
		16#28f4# => X"e3120510",
		16#28f5# => X"130dc10f",
		16#28f6# => X"8327c10b",
		16#28f7# => X"63c64701",
		16#28f8# => X"93771400",
		16#28f9# => X"63820722",
		16#28fa# => X"83278103",
		16#28fb# => X"03274102",
		16#28fc# => X"130d8d00",
		16#28fd# => X"232cfdfe",
		16#28fe# => X"83274102",
		16#28ff# => X"232efdfe",
		16#2900# => X"8327c10d",
		16#2901# => X"b387e700",
		16#2902# => X"232ef10c",
		16#2903# => X"8327810d",
		16#2904# => X"13077000",
		16#2905# => X"93871700",
		16#2906# => X"232cf10c",
		16#2907# => X"635ef700",
		16#2908# => X"1306410d",
		16#2909# => X"93850900",
		16#290a# => X"13050900",
		16#290b# => X"ef105061",
		16#290c# => X"e312050a",
		16#290d# => X"130dc10f",
		16#290e# => X"9304faff",
		16#290f# => X"6356901c",
		16#2910# => X"930a0001",
		16#2911# => X"930b7000",
		16#2912# => X"03268101",
		16#2913# => X"8327810d",
		16#2914# => X"0327c10d",
		16#2915# => X"2320cd00",
		16#2916# => X"93871700",
		16#2917# => X"93068d00",
		16#2918# => X"63c29a02",
		16#2919# => X"23229d00",
		16#291a# => X"b384e400",
		16#291b# => X"232e910c",
		16#291c# => X"232cf10c",
		16#291d# => X"13077000",
		16#291e# => X"138d0600",
		16#291f# => X"6356f718",
		16#2920# => X"6fe09fff",
		16#2921# => X"13070701",
		16#2922# => X"23225d01",
		16#2923# => X"232ee10c",
		16#2924# => X"232cf10c",
		16#2925# => X"63defb00",
		16#2926# => X"1306410d",
		16#2927# => X"93850900",
		16#2928# => X"13050900",
		16#2929# => X"ef10d059",
		16#292a# => X"e3160502",
		16#292b# => X"9306c10f",
		16#292c# => X"938404ff",
		16#292d# => X"138d0600",
		16#292e# => X"6ff01ff9",
		16#292f# => X"0327c10b",
		16#2930# => X"634ae01c",
		16#2931# => X"b7470110",
		16#2932# => X"9387c792",
		16#2933# => X"2320fd00",
		16#2934# => X"93071000",
		16#2935# => X"2322fd00",
		16#2936# => X"8327810d",
		16#2937# => X"938d1d00",
		16#2938# => X"232eb10d",
		16#2939# => X"93871700",
		16#293a# => X"232cf10c",
		16#293b# => X"13077000",
		16#293c# => X"130d8d00",
		16#293d# => X"635ef700",
		16#293e# => X"1306410d",
		16#293f# => X"93850900",
		16#2940# => X"13050900",
		16#2941# => X"ef10d053",
		16#2942# => X"6316057c",
		16#2943# => X"130dc10f",
		16#2944# => X"8327c10b",
		16#2945# => X"63980700",
		16#2946# => X"63160a00",
		16#2947# => X"93771400",
		16#2948# => X"6384070e",
		16#2949# => X"83278103",
		16#294a# => X"03274102",
		16#294b# => X"93088d00",
		16#294c# => X"2320fd00",
		16#294d# => X"83274102",
		16#294e# => X"2322fd00",
		16#294f# => X"8327c10d",
		16#2950# => X"b387e700",
		16#2951# => X"232ef10c",
		16#2952# => X"8327810d",
		16#2953# => X"13077000",
		16#2954# => X"93871700",
		16#2955# => X"232cf10c",
		16#2956# => X"635ef700",
		16#2957# => X"1306410d",
		16#2958# => X"93850900",
		16#2959# => X"13050900",
		16#295a# => X"ef10904d",
		16#295b# => X"63140576",
		16#295c# => X"9308c10f",
		16#295d# => X"832ac10b",
		16#295e# => X"63d00a06",
		16#295f# => X"b30a5041",
		16#2960# => X"13870800",
		16#2961# => X"930b0001",
		16#2962# => X"130c7000",
		16#2963# => X"03268101",
		16#2964# => X"8327810d",
		16#2965# => X"8326c10d",
		16#2966# => X"2320c700",
		16#2967# => X"93871700",
		16#2968# => X"93888800",
		16#2969# => X"63cc5b0b",
		16#296a# => X"23225701",
		16#296b# => X"b38ada00",
		16#296c# => X"232e510d",
		16#296d# => X"232cf10c",
		16#296e# => X"13077000",
		16#296f# => X"635ef700",
		16#2970# => X"1306410d",
		16#2971# => X"93850900",
		16#2972# => X"13050900",
		16#2973# => X"ef105047",
		16#2974# => X"63120570",
		16#2975# => X"9308c10f",
		16#2976# => X"8327c10d",
		16#2977# => X"23a09800",
		16#2978# => X"23a24801",
		16#2979# => X"b3874701",
		16#297a# => X"232ef10c",
		16#297b# => X"8327810d",
		16#297c# => X"13077000",
		16#297d# => X"138d8800",
		16#297e# => X"93871700",
		16#297f# => X"232cf10c",
		16#2980# => X"6354f700",
		16#2981# => X"6fe05fe7",
		16#2982# => X"13744400",
		16#2983# => X"63140466",
		16#2984# => X"032dc102",
		16#2985# => X"83270103",
		16#2986# => X"6354fd00",
		16#2987# => X"138d0700",
		16#2988# => X"83278102",
		16#2989# => X"b387a701",
		16#298a# => X"2324f102",
		16#298b# => X"8327c10d",
		16#298c# => X"638c0700",
		16#298d# => X"1306410d",
		16#298e# => X"93850900",
		16#298f# => X"13050900",
		16#2990# => X"ef101040",
		16#2991# => X"63180568",
		16#2992# => X"83270101",
		16#2993# => X"232c010c",
		16#2994# => X"639c076c",
		16#2995# => X"130dc10f",
		16#2996# => X"6ff01f84",
		16#2997# => X"93860601",
		16#2998# => X"23227701",
		16#2999# => X"232ed10c",
		16#299a# => X"232cf10c",
		16#299b# => X"635efc00",
		16#299c# => X"1306410d",
		16#299d# => X"93850900",
		16#299e# => X"13050900",
		16#299f# => X"ef10503c",
		16#29a0# => X"631a0564",
		16#29a1# => X"9308c10f",
		16#29a2# => X"938a0aff",
		16#29a3# => X"13870800",
		16#29a4# => X"6ff0dfef",
		16#29a5# => X"938a0c00",
		16#29a6# => X"63549a01",
		16#29a7# => X"930a0a00",
		16#29a8# => X"63525005",
		16#29a9# => X"0327810d",
		16#29aa# => X"b38dba01",
		16#29ab# => X"23209d00",
		16#29ac# => X"13071700",
		16#29ad# => X"23225d01",
		16#29ae# => X"232eb10d",
		16#29af# => X"232ce10c",
		16#29b0# => X"93067000",
		16#29b1# => X"130d8d00",
		16#29b2# => X"63dee600",
		16#29b3# => X"1306410d",
		16#29b4# => X"93850900",
		16#29b5# => X"13050900",
		16#29b6# => X"ef109036",
		16#29b7# => X"631c055e",
		16#29b8# => X"130dc10f",
		16#29b9# => X"63d40a00",
		16#29ba# => X"930a0000",
		16#29bb# => X"b38a5c41",
		16#29bc# => X"635e5005",
		16#29bd# => X"130b0001",
		16#29be# => X"930d7000",
		16#29bf# => X"83278101",
		16#29c0# => X"0327810d",
		16#29c1# => X"8326c10d",
		16#29c2# => X"2320fd00",
		16#29c3# => X"13071700",
		16#29c4# => X"13068d00",
		16#29c5# => X"634c5b19",
		16#29c6# => X"23225d01",
		16#29c7# => X"b38ada00",
		16#29c8# => X"232e510d",
		16#29c9# => X"232ce10c",
		16#29ca# => X"93067000",
		16#29cb# => X"130d0600",
		16#29cc# => X"63dee600",
		16#29cd# => X"1306410d",
		16#29ce# => X"93850900",
		16#29cf# => X"13050900",
		16#29d0# => X"ef101030",
		16#29d1# => X"63180558",
		16#29d2# => X"130dc10f",
		16#29d3# => X"93770440",
		16#29d4# => X"b38a9401",
		16#29d5# => X"63800702",
		16#29d6# => X"130b7000",
		16#29d7# => X"b38d4401",
		16#29d8# => X"63920b18",
		16#29d9# => X"63120c18",
		16#29da# => X"b3874401",
		16#29db# => X"63f45701",
		16#29dc# => X"938a0700",
		16#29dd# => X"8327c10b",
		16#29de# => X"63c64701",
		16#29df# => X"93771400",
		16#29e0# => X"638a0704",
		16#29e1# => X"83278103",
		16#29e2# => X"03274102",
		16#29e3# => X"130d8d00",
		16#29e4# => X"232cfdfe",
		16#29e5# => X"83274102",
		16#29e6# => X"232efdfe",
		16#29e7# => X"8327c10d",
		16#29e8# => X"b387e700",
		16#29e9# => X"232ef10c",
		16#29ea# => X"8327810d",
		16#29eb# => X"13077000",
		16#29ec# => X"93871700",
		16#29ed# => X"232cf10c",
		16#29ee# => X"635ef700",
		16#29ef# => X"1306410d",
		16#29f0# => X"93850900",
		16#29f1# => X"13050900",
		16#29f2# => X"ef109027",
		16#29f3# => X"63140550",
		16#29f4# => X"130dc10f",
		16#29f5# => X"b3844401",
		16#29f6# => X"b3875441",
		16#29f7# => X"8324c10b",
		16#29f8# => X"b3049a40",
		16#29f9# => X"63d49700",
		16#29fa# => X"93840700",
		16#29fb# => X"63549004",
		16#29fc# => X"8327c10d",
		16#29fd# => X"23205d01",
		16#29fe# => X"23229d00",
		16#29ff# => X"b387f400",
		16#2a00# => X"232ef10c",
		16#2a01# => X"8327810d",
		16#2a02# => X"13077000",
		16#2a03# => X"130d8d00",
		16#2a04# => X"93871700",
		16#2a05# => X"232cf10c",
		16#2a06# => X"635ef700",
		16#2a07# => X"1306410d",
		16#2a08# => X"93850900",
		16#2a09# => X"13050900",
		16#2a0a# => X"ef109021",
		16#2a0b# => X"6314054a",
		16#2a0c# => X"130dc10f",
		16#2a0d# => X"93870400",
		16#2a0e# => X"63d40400",
		16#2a0f# => X"93070000",
		16#2a10# => X"8324c10b",
		16#2a11# => X"b3049a40",
		16#2a12# => X"b384f440",
		16#2a13# => X"e35e90da",
		16#2a14# => X"930a0001",
		16#2a15# => X"930b7000",
		16#2a16# => X"03268101",
		16#2a17# => X"8327810d",
		16#2a18# => X"0327c10d",
		16#2a19# => X"2320cd00",
		16#2a1a# => X"93871700",
		16#2a1b# => X"93068d00",
		16#2a1c# => X"e3da9abe",
		16#2a1d# => X"13070701",
		16#2a1e# => X"23225d01",
		16#2a1f# => X"232ee10c",
		16#2a20# => X"232cf10c",
		16#2a21# => X"63defb00",
		16#2a22# => X"1306410d",
		16#2a23# => X"93850900",
		16#2a24# => X"13050900",
		16#2a25# => X"ef10d01a",
		16#2a26# => X"631e0542",
		16#2a27# => X"9306c10f",
		16#2a28# => X"938404ff",
		16#2a29# => X"138d0600",
		16#2a2a# => X"6ff01ffb",
		16#2a2b# => X"93860601",
		16#2a2c# => X"23226d01",
		16#2a2d# => X"232ed10c",
		16#2a2e# => X"232ce10c",
		16#2a2f# => X"63deed00",
		16#2a30# => X"1306410d",
		16#2a31# => X"93850900",
		16#2a32# => X"13050900",
		16#2a33# => X"ef105017",
		16#2a34# => X"63120540",
		16#2a35# => X"1306c10f",
		16#2a36# => X"938a0aff",
		16#2a37# => X"130d0600",
		16#2a38# => X"6ff0dfe1",
		16#2a39# => X"63020c0e",
		16#2a3a# => X"130cfcff",
		16#2a3b# => X"8327c103",
		16#2a3c# => X"03274103",
		16#2a3d# => X"130d8d00",
		16#2a3e# => X"232cfdfe",
		16#2a3f# => X"83274103",
		16#2a40# => X"232efdfe",
		16#2a41# => X"8327c10d",
		16#2a42# => X"b387e700",
		16#2a43# => X"232ef10c",
		16#2a44# => X"8327810d",
		16#2a45# => X"93871700",
		16#2a46# => X"232cf10c",
		16#2a47# => X"635efb00",
		16#2a48# => X"1306410d",
		16#2a49# => X"93850900",
		16#2a4a# => X"13050900",
		16#2a4b# => X"ef105011",
		16#2a4c# => X"6312053a",
		16#2a4d# => X"130dc10f",
		16#2a4e# => X"83274101",
		16#2a4f# => X"33875d41",
		16#2a50# => X"83c70700",
		16#2a51# => X"6354f700",
		16#2a52# => X"93070700",
		16#2a53# => X"6356f004",
		16#2a54# => X"0327c10d",
		16#2a55# => X"23205d01",
		16#2a56# => X"2322fd00",
		16#2a57# => X"3387e700",
		16#2a58# => X"232ee10c",
		16#2a59# => X"0327810d",
		16#2a5a# => X"130d8d00",
		16#2a5b# => X"13071700",
		16#2a5c# => X"232ce10c",
		16#2a5d# => X"6352eb02",
		16#2a5e# => X"1306410d",
		16#2a5f# => X"93850900",
		16#2a60# => X"13050900",
		16#2a61# => X"2326f100",
		16#2a62# => X"ef10900b",
		16#2a63# => X"63140534",
		16#2a64# => X"8327c100",
		16#2a65# => X"130dc10f",
		16#2a66# => X"13870700",
		16#2a67# => X"63d40700",
		16#2a68# => X"13070000",
		16#2a69# => X"83274101",
		16#2a6a# => X"13080001",
		16#2a6b# => X"83c70700",
		16#2a6c# => X"b387e740",
		16#2a6d# => X"6346f006",
		16#2a6e# => X"83274101",
		16#2a6f# => X"83c70700",
		16#2a70# => X"b38afa00",
		16#2a71# => X"6ff0dfd9",
		16#2a72# => X"83274101",
		16#2a73# => X"938bfbff",
		16#2a74# => X"9387f7ff",
		16#2a75# => X"232af100",
		16#2a76# => X"6ff05ff1",
		16#2a77# => X"93860601",
		16#2a78# => X"23220d01",
		16#2a79# => X"232ed10c",
		16#2a7a# => X"232ce10c",
		16#2a7b# => X"6356eb02",
		16#2a7c# => X"1306410d",
		16#2a7d# => X"93850900",
		16#2a7e# => X"13050900",
		16#2a7f# => X"23240105",
		16#2a80# => X"2326f100",
		16#2a81# => X"ef10d003",
		16#2a82# => X"6316052c",
		16#2a83# => X"03288104",
		16#2a84# => X"8327c100",
		16#2a85# => X"1306c10f",
		16#2a86# => X"938707ff",
		16#2a87# => X"130d0600",
		16#2a88# => X"83258101",
		16#2a89# => X"0327810d",
		16#2a8a# => X"8326c10d",
		16#2a8b# => X"2320bd00",
		16#2a8c# => X"13071700",
		16#2a8d# => X"13068d00",
		16#2a8e# => X"e342f8fa",
		16#2a8f# => X"2322fd00",
		16#2a90# => X"b387d700",
		16#2a91# => X"232ef10c",
		16#2a92# => X"232ce10c",
		16#2a93# => X"130d0600",
		16#2a94# => X"e354ebf6",
		16#2a95# => X"1306410d",
		16#2a96# => X"93850900",
		16#2a97# => X"13050900",
		16#2a98# => X"ef10007e",
		16#2a99# => X"63180526",
		16#2a9a# => X"130dc10f",
		16#2a9b# => X"6ff0dff4",
		16#2a9c# => X"8327810d",
		16#2a9d# => X"13071000",
		16#2a9e# => X"23209d00",
		16#2a9f# => X"938d1d00",
		16#2aa0# => X"93871700",
		16#2aa1# => X"930b8d00",
		16#2aa2# => X"63464701",
		16#2aa3# => X"93761400",
		16#2aa4# => X"6386061c",
		16#2aa5# => X"13071000",
		16#2aa6# => X"2322ed00",
		16#2aa7# => X"232eb10d",
		16#2aa8# => X"232cf10c",
		16#2aa9# => X"13077000",
		16#2aaa# => X"635ef700",
		16#2aab# => X"1306410d",
		16#2aac# => X"93850900",
		16#2aad# => X"13050900",
		16#2aae# => X"ef108078",
		16#2aaf# => X"631c0520",
		16#2ab0# => X"930bc10f",
		16#2ab1# => X"83278103",
		16#2ab2# => X"03274102",
		16#2ab3# => X"938b8b00",
		16#2ab4# => X"23acfbfe",
		16#2ab5# => X"83274102",
		16#2ab6# => X"23aefbfe",
		16#2ab7# => X"8327c10d",
		16#2ab8# => X"b387e700",
		16#2ab9# => X"232ef10c",
		16#2aba# => X"8327810d",
		16#2abb# => X"13077000",
		16#2abc# => X"93871700",
		16#2abd# => X"232cf10c",
		16#2abe# => X"635ef700",
		16#2abf# => X"1306410d",
		16#2ac0# => X"93850900",
		16#2ac1# => X"13050900",
		16#2ac2# => X"ef108073",
		16#2ac3# => X"6314051c",
		16#2ac4# => X"930bc10f",
		16#2ac5# => X"8327010e",
		16#2ac6# => X"93050109",
		16#2ac7# => X"1305010a",
		16#2ac8# => X"2320f10a",
		16#2ac9# => X"8327410e",
		16#2aca# => X"930afaff",
		16#2acb# => X"23280108",
		16#2acc# => X"2322f10a",
		16#2acd# => X"8327810e",
		16#2ace# => X"232a0108",
		16#2acf# => X"232c0108",
		16#2ad0# => X"2324f10a",
		16#2ad1# => X"8327c10e",
		16#2ad2# => X"232e0108",
		16#2ad3# => X"2326f10a",
		16#2ad4# => X"ef408056",
		16#2ad5# => X"63060508",
		16#2ad6# => X"8327c10d",
		16#2ad7# => X"0327810d",
		16#2ad8# => X"93841400",
		16#2ad9# => X"9387f7ff",
		16#2ada# => X"b3874701",
		16#2adb# => X"13071700",
		16#2adc# => X"23a09b00",
		16#2add# => X"23a25b01",
		16#2ade# => X"232ef10c",
		16#2adf# => X"232ce10c",
		16#2ae0# => X"93077000",
		16#2ae1# => X"938b8b00",
		16#2ae2# => X"63dee700",
		16#2ae3# => X"1306410d",
		16#2ae4# => X"93850900",
		16#2ae5# => X"13050900",
		16#2ae6# => X"ef10806a",
		16#2ae7# => X"631c0512",
		16#2ae8# => X"930bc10f",
		16#2ae9# => X"9307410c",
		16#2aea# => X"23a0fb00",
		16#2aeb# => X"83270104",
		16#2aec# => X"03270104",
		16#2aed# => X"138d8b00",
		16#2aee# => X"23a2fb00",
		16#2aef# => X"8327c10d",
		16#2af0# => X"b387e700",
		16#2af1# => X"232ef10c",
		16#2af2# => X"8327810d",
		16#2af3# => X"13077000",
		16#2af4# => X"93871700",
		16#2af5# => X"232cf10c",
		16#2af6# => X"e358f7a2",
		16#2af7# => X"6fe0df89",
		16#2af8# => X"e35250fd",
		16#2af9# => X"93040001",
		16#2afa# => X"130c7000",
		16#2afb# => X"03268101",
		16#2afc# => X"0327810d",
		16#2afd# => X"8327c10d",
		16#2afe# => X"23a0cb00",
		16#2aff# => X"13071700",
		16#2b00# => X"93868b00",
		16#2b01# => X"63c05403",
		16#2b02# => X"b387fa00",
		16#2b03# => X"23a25b01",
		16#2b04# => X"232ef10c",
		16#2b05# => X"232ce10c",
		16#2b06# => X"93077000",
		16#2b07# => X"938b0600",
		16#2b08# => X"6ff09ff6",
		16#2b09# => X"93870701",
		16#2b0a# => X"23a29b00",
		16#2b0b# => X"232ef10c",
		16#2b0c# => X"232ce10c",
		16#2b0d# => X"635eec00",
		16#2b0e# => X"1306410d",
		16#2b0f# => X"93850900",
		16#2b10# => X"13050900",
		16#2b11# => X"ef10c05f",
		16#2b12# => X"63160508",
		16#2b13# => X"9306c10f",
		16#2b14# => X"938a0aff",
		16#2b15# => X"938b0600",
		16#2b16# => X"6ff05ff9",
		16#2b17# => X"2322ed00",
		16#2b18# => X"232eb10d",
		16#2b19# => X"232cf10c",
		16#2b1a# => X"13077000",
		16#2b1b# => X"e35cf7f2",
		16#2b1c# => X"6ff0dff1",
		16#2b1d# => X"8327c102",
		16#2b1e# => X"03270103",
		16#2b1f# => X"3384e740",
		16#2b20# => X"e3588098",
		16#2b21# => X"b7440110",
		16#2b22# => X"930a0001",
		16#2b23# => X"9384c41c",
		16#2b24# => X"930b7000",
		16#2b25# => X"8327810d",
		16#2b26# => X"23209d00",
		16#2b27# => X"0327c10d",
		16#2b28# => X"93871700",
		16#2b29# => X"63c68a04",
		16#2b2a# => X"23228d00",
		16#2b2b# => X"3304e400",
		16#2b2c# => X"232e810c",
		16#2b2d# => X"232cf10c",
		16#2b2e# => X"13077000",
		16#2b2f# => X"e35af794",
		16#2b30# => X"1306410d",
		16#2b31# => X"93850900",
		16#2b32# => X"13050900",
		16#2b33# => X"ef104057",
		16#2b34# => X"e3000594",
		16#2b35# => X"83270101",
		16#2b36# => X"63940700",
		16#2b37# => X"6fe05fa0",
		16#2b38# => X"93850700",
		16#2b39# => X"13050900",
		16#2b3a# => X"ef904fcb",
		16#2b3b# => X"6fe05f9f",
		16#2b3c# => X"13070701",
		16#2b3d# => X"23225d01",
		16#2b3e# => X"232ee10c",
		16#2b3f# => X"232cf10c",
		16#2b40# => X"130d8d00",
		16#2b41# => X"63defb00",
		16#2b42# => X"1306410d",
		16#2b43# => X"93850900",
		16#2b44# => X"13050900",
		16#2b45# => X"ef10c052",
		16#2b46# => X"e31e05fa",
		16#2b47# => X"130dc10f",
		16#2b48# => X"130404ff",
		16#2b49# => X"6ff01ff7",
		16#2b4a# => X"83250101",
		16#2b4b# => X"13050900",
		16#2b4c# => X"ef90cfc6",
		16#2b4d# => X"6ff01f92",
		16#2b4e# => X"8327c10d",
		16#2b4f# => X"63940700",
		16#2b50# => X"6fe01f9a",
		16#2b51# => X"1306410d",
		16#2b52# => X"93850900",
		16#2b53# => X"13050900",
		16#2b54# => X"ef10004f",
		16#2b55# => X"6fe0df98",
		16#2b56# => X"83278600",
		16#2b57# => X"130101fd",
		16#2b58# => X"23248102",
		16#2b59# => X"23261102",
		16#2b5a# => X"23229102",
		16#2b5b# => X"23202103",
		16#2b5c# => X"232e3101",
		16#2b5d# => X"232c4101",
		16#2b5e# => X"232a5101",
		16#2b5f# => X"23286101",
		16#2b60# => X"23267101",
		16#2b61# => X"23248101",
		16#2b62# => X"13040600",
		16#2b63# => X"639e0702",
		16#2b64# => X"23220600",
		16#2b65# => X"13050000",
		16#2b66# => X"8320c102",
		16#2b67# => X"03248102",
		16#2b68# => X"83244102",
		16#2b69# => X"03290102",
		16#2b6a# => X"8329c101",
		16#2b6b# => X"032a8101",
		16#2b6c# => X"832a4101",
		16#2b6d# => X"032b0101",
		16#2b6e# => X"832bc100",
		16#2b6f# => X"032c8100",
		16#2b70# => X"13010103",
		16#2b71# => X"67800000",
		16#2b72# => X"83a74506",
		16#2b73# => X"13890500",
		16#2b74# => X"13972701",
		16#2b75# => X"635a0706",
		16#2b76# => X"83240600",
		16#2b77# => X"130a0500",
		16#2b78# => X"930bf0ff",
		16#2b79# => X"83278400",
		16#2b7a# => X"639a0700",
		16#2b7b# => X"13050000",
		16#2b7c# => X"23240400",
		16#2b7d# => X"23220400",
		16#2b7e# => X"6ff01ffa",
		16#2b7f# => X"83a94400",
		16#2b80# => X"03ab0400",
		16#2b81# => X"930a0000",
		16#2b82# => X"13dc2900",
		16#2b83# => X"63ce8a01",
		16#2b84# => X"83278400",
		16#2b85# => X"93f9c9ff",
		16#2b86# => X"93848400",
		16#2b87# => X"b3893741",
		16#2b88# => X"23243401",
		16#2b89# => X"6ff01ffc",
		16#2b8a# => X"83250b00",
		16#2b8b# => X"13060900",
		16#2b8c# => X"13050a00",
		16#2b8d# => X"ef10c00f",
		16#2b8e# => X"130b4b00",
		16#2b8f# => X"630a7501",
		16#2b90# => X"938a1a00",
		16#2b91# => X"6ff09ffc",
		16#2b92# => X"ef900fdb",
		16#2b93# => X"6ff05ffa",
		16#2b94# => X"1305f0ff",
		16#2b95# => X"6ff0dff9",
		16#2b96# => X"130101ed",
		16#2b97# => X"23248112",
		16#2b98# => X"232e3111",
		16#2b99# => X"232c4111",
		16#2b9a# => X"2320a111",
		16#2b9b# => X"23261112",
		16#2b9c# => X"23229112",
		16#2b9d# => X"23202113",
		16#2b9e# => X"232a5111",
		16#2b9f# => X"23286111",
		16#2ba0# => X"23267111",
		16#2ba1# => X"23248111",
		16#2ba2# => X"23229111",
		16#2ba3# => X"232eb10f",
		16#2ba4# => X"93090500",
		16#2ba5# => X"13840500",
		16#2ba6# => X"130a0600",
		16#2ba7# => X"138d0600",
		16#2ba8# => X"63080500",
		16#2ba9# => X"83278503",
		16#2baa# => X"63940700",
		16#2bab# => X"ef90cf83",
		16#2bac# => X"8317c400",
		16#2bad# => X"13972701",
		16#2bae# => X"63420702",
		16#2baf# => X"b7260000",
		16#2bb0# => X"03274406",
		16#2bb1# => X"b3e7d700",
		16#2bb2# => X"2316f400",
		16#2bb3# => X"b7e7ffff",
		16#2bb4# => X"9387f7ff",
		16#2bb5# => X"b377f700",
		16#2bb6# => X"2322f406",
		16#2bb7# => X"8357c400",
		16#2bb8# => X"93f78700",
		16#2bb9# => X"638e0706",
		16#2bba# => X"83270401",
		16#2bbb# => X"638a0706",
		16#2bbc# => X"8357c400",
		16#2bbd# => X"1307a000",
		16#2bbe# => X"93f7a701",
		16#2bbf# => X"6390e708",
		16#2bc0# => X"8317e400",
		16#2bc1# => X"63cc0706",
		16#2bc2# => X"93060d00",
		16#2bc3# => X"13060a00",
		16#2bc4# => X"93050400",
		16#2bc5# => X"13850900",
		16#2bc6# => X"ef00503c",
		16#2bc7# => X"2320a100",
		16#2bc8# => X"8320c112",
		16#2bc9# => X"03248112",
		16#2bca# => X"03250100",
		16#2bcb# => X"83244112",
		16#2bcc# => X"03290112",
		16#2bcd# => X"8329c111",
		16#2bce# => X"032a8111",
		16#2bcf# => X"832a4111",
		16#2bd0# => X"032b0111",
		16#2bd1# => X"832bc110",
		16#2bd2# => X"032c8110",
		16#2bd3# => X"832c4110",
		16#2bd4# => X"032d0110",
		16#2bd5# => X"832dc10f",
		16#2bd6# => X"13010113",
		16#2bd7# => X"67800000",
		16#2bd8# => X"93050400",
		16#2bd9# => X"13850900",
		16#2bda# => X"ef809faa",
		16#2bdb# => X"e30205f8",
		16#2bdc# => X"9307f0ff",
		16#2bdd# => X"2320f100",
		16#2bde# => X"6ff09ffa",
		16#2bdf# => X"9307c104",
		16#2be0# => X"2320f104",
		16#2be1# => X"938b0700",
		16#2be2# => X"b7470110",
		16#2be3# => X"9387c71e",
		16#2be4# => X"232ef100",
		16#2be5# => X"b7470110",
		16#2be6# => X"93878736",
		16#2be7# => X"23240104",
		16#2be8# => X"23220104",
		16#2be9# => X"23240100",
		16#2bea# => X"23220100",
		16#2beb# => X"23260100",
		16#2bec# => X"232a0100",
		16#2bed# => X"23200100",
		16#2bee# => X"2328f100",
		16#2bef# => X"93040a00",
		16#2bf0# => X"93065002",
		16#2bf1# => X"83c70400",
		16#2bf2# => X"63840700",
		16#2bf3# => X"6392d70a",
		16#2bf4# => X"33894441",
		16#2bf5# => X"630a0904",
		16#2bf6# => X"83278104",
		16#2bf7# => X"23a04b01",
		16#2bf8# => X"23a22b01",
		16#2bf9# => X"b3872701",
		16#2bfa# => X"2324f104",
		16#2bfb# => X"83274104",
		16#2bfc# => X"93067000",
		16#2bfd# => X"938b8b00",
		16#2bfe# => X"93871700",
		16#2bff# => X"2322f104",
		16#2c00# => X"63def600",
		16#2c01# => X"13060104",
		16#2c02# => X"93050400",
		16#2c03# => X"13850900",
		16#2c04# => X"eff09fd4",
		16#2c05# => X"e3180524",
		16#2c06# => X"930bc104",
		16#2c07# => X"83270100",
		16#2c08# => X"b3872701",
		16#2c09# => X"2320f100",
		16#2c0a# => X"83c70400",
		16#2c0b# => X"e3800728",
		16#2c0c# => X"138a1400",
		16#2c0d# => X"a30d0102",
		16#2c0e# => X"1309f0ff",
		16#2c0f# => X"930a0000",
		16#2c10# => X"130b0000",
		16#2c11# => X"93049000",
		16#2c12# => X"930ca005",
		16#2c13# => X"834d0a00",
		16#2c14# => X"130a1a00",
		16#2c15# => X"93860dfe",
		16#2c16# => X"e3e0dc0c",
		16#2c17# => X"8327c101",
		16#2c18# => X"93962600",
		16#2c19# => X"b386f600",
		16#2c1a# => X"83a60600",
		16#2c1b# => X"67800600",
		16#2c1c# => X"93841400",
		16#2c1d# => X"6ff01ff5",
		16#2c1e# => X"b7460110",
		16#2c1f# => X"93878691",
		16#2c20# => X"2324f100",
		16#2c21# => X"93760b02",
		16#2c22# => X"638e066a",
		16#2c23# => X"130d7d00",
		16#2c24# => X"137d8dff",
		16#2c25# => X"83280d00",
		16#2c26# => X"832c4d00",
		16#2c27# => X"130c8d00",
		16#2c28# => X"93761b00",
		16#2c29# => X"638e0600",
		16#2c2a# => X"b3e69801",
		16#2c2b# => X"638a0600",
		16#2c2c# => X"93060003",
		16#2c2d# => X"230ed102",
		16#2c2e# => X"a30eb103",
		16#2c2f# => X"136b2b00",
		16#2c30# => X"137bfbbf",
		16#2c31# => X"6f008033",
		16#2c32# => X"13850900",
		16#2c33# => X"efb05f96",
		16#2c34# => X"83274500",
		16#2c35# => X"13850700",
		16#2c36# => X"232af100",
		16#2c37# => X"ef608ff3",
		16#2c38# => X"2326a100",
		16#2c39# => X"13850900",
		16#2c3a# => X"efb09f94",
		16#2c3b# => X"83278500",
		16#2c3c# => X"2322f100",
		16#2c3d# => X"8327c100",
		16#2c3e# => X"e38807f4",
		16#2c3f# => X"83274100",
		16#2c40# => X"e38407f4",
		16#2c41# => X"83c60700",
		16#2c42# => X"e38006f4",
		16#2c43# => X"136b0b40",
		16#2c44# => X"6ff09ff3",
		16#2c45# => X"8346b103",
		16#2c46# => X"e39806f2",
		16#2c47# => X"93060002",
		16#2c48# => X"a30dd102",
		16#2c49# => X"6ff05ff2",
		16#2c4a# => X"136b1b00",
		16#2c4b# => X"6ff0dff1",
		16#2c4c# => X"832a0d00",
		16#2c4d# => X"130d4d00",
		16#2c4e# => X"e3d80af0",
		16#2c4f# => X"b30a5041",
		16#2c50# => X"136b4b00",
		16#2c51# => X"6ff05ff0",
		16#2c52# => X"9306b002",
		16#2c53# => X"6ff05ffd",
		16#2c54# => X"834d0a00",
		16#2c55# => X"9307a002",
		16#2c56# => X"130c1a00",
		16#2c57# => X"6394fd04",
		16#2c58# => X"03290d00",
		16#2c59# => X"13064d00",
		16#2c5a# => X"63540900",
		16#2c5b# => X"1309f0ff",
		16#2c5c# => X"130d0600",
		16#2c5d# => X"130a0c00",
		16#2c5e# => X"6ff01fed",
		16#2c5f# => X"13050900",
		16#2c60# => X"9305a000",
		16#2c61# => X"130c1c00",
		16#2c62# => X"ef70804a",
		16#2c63# => X"834dfcff",
		16#2c64# => X"33094501",
		16#2c65# => X"138a0dfd",
		16#2c66# => X"e3f244ff",
		16#2c67# => X"130a0c00",
		16#2c68# => X"6ff05feb",
		16#2c69# => X"13090000",
		16#2c6a# => X"6ff0dffe",
		16#2c6b# => X"136b0b08",
		16#2c6c# => X"6ff09fe9",
		16#2c6d# => X"130c0a00",
		16#2c6e# => X"930a0000",
		16#2c6f# => X"13850a00",
		16#2c70# => X"9305a000",
		16#2c71# => X"130c1c00",
		16#2c72# => X"ef708046",
		16#2c73# => X"938a0dfd",
		16#2c74# => X"834dfcff",
		16#2c75# => X"b38aaa00",
		16#2c76# => X"13860dfd",
		16#2c77# => X"e3f0c4fe",
		16#2c78# => X"6ff0dffb",
		16#2c79# => X"03460a00",
		16#2c7a# => X"93068006",
		16#2c7b# => X"6318d600",
		16#2c7c# => X"130a1a00",
		16#2c7d# => X"136b0b20",
		16#2c7e# => X"6ff01fe5",
		16#2c7f# => X"136b0b04",
		16#2c80# => X"6ff09fe4",
		16#2c81# => X"03460a00",
		16#2c82# => X"9306c006",
		16#2c83# => X"6318d600",
		16#2c84# => X"130a1a00",
		16#2c85# => X"136b0b02",
		16#2c86# => X"6ff01fe3",
		16#2c87# => X"136b0b01",
		16#2c88# => X"6ff09fe2",
		16#2c89# => X"83260d00",
		16#2c8a# => X"130c4d00",
		16#2c8b# => X"a30d0102",
		16#2c8c# => X"2306d108",
		16#2c8d# => X"13091000",
		16#2c8e# => X"930c0000",
		16#2c8f# => X"9304c108",
		16#2c90# => X"6f00401f",
		16#2c91# => X"136b0b01",
		16#2c92# => X"93760b02",
		16#2c93# => X"638c0604",
		16#2c94# => X"130d7d00",
		16#2c95# => X"137d8dff",
		16#2c96# => X"83280d00",
		16#2c97# => X"832c4d00",
		16#2c98# => X"130c8d00",
		16#2c99# => X"63de0c00",
		16#2c9a# => X"b3081041",
		16#2c9b# => X"b3361001",
		16#2c9c# => X"33039041",
		16#2c9d# => X"b30cd340",
		16#2c9e# => X"9306d002",
		16#2c9f# => X"a30dd102",
		16#2ca0# => X"9306f0ff",
		16#2ca1# => X"631cd94e",
		16#2ca2# => X"63960c56",
		16#2ca3# => X"93069000",
		16#2ca4# => X"63e21657",
		16#2ca5# => X"93880803",
		16#2ca6# => X"a307110f",
		16#2ca7# => X"9304f10e",
		16#2ca8# => X"6f00c053",
		16#2ca9# => X"93760b01",
		16#2caa# => X"130c4d00",
		16#2cab# => X"63880600",
		16#2cac# => X"83280d00",
		16#2cad# => X"93dcf841",
		16#2cae# => X"6ff0dffa",
		16#2caf# => X"93760b04",
		16#2cb0# => X"83280d00",
		16#2cb1# => X"63880600",
		16#2cb2# => X"93980801",
		16#2cb3# => X"93d80841",
		16#2cb4# => X"6ff05ffe",
		16#2cb5# => X"93760b20",
		16#2cb6# => X"e38e06fc",
		16#2cb7# => X"93988801",
		16#2cb8# => X"93d88841",
		16#2cb9# => X"6ff01ffd",
		16#2cba# => X"13760b02",
		16#2cbb# => X"83260d00",
		16#2cbc# => X"130d4d00",
		16#2cbd# => X"630c0600",
		16#2cbe# => X"83270100",
		16#2cbf# => X"23a0f600",
		16#2cc0# => X"93d7f741",
		16#2cc1# => X"23a2f600",
		16#2cc2# => X"6ff05fcb",
		16#2cc3# => X"13760b01",
		16#2cc4# => X"63080600",
		16#2cc5# => X"83270100",
		16#2cc6# => X"23a0f600",
		16#2cc7# => X"6ff01fca",
		16#2cc8# => X"13760b04",
		16#2cc9# => X"63080600",
		16#2cca# => X"83570100",
		16#2ccb# => X"2390f600",
		16#2ccc# => X"6ff0dfc8",
		16#2ccd# => X"93770b20",
		16#2cce# => X"e38e07fc",
		16#2ccf# => X"83470100",
		16#2cd0# => X"2380f600",
		16#2cd1# => X"6ff09fc7",
		16#2cd2# => X"136b0b01",
		16#2cd3# => X"93760b02",
		16#2cd4# => X"63860604",
		16#2cd5# => X"130d7d00",
		16#2cd6# => X"137d8dff",
		16#2cd7# => X"83280d00",
		16#2cd8# => X"832c4d00",
		16#2cd9# => X"130c8d00",
		16#2cda# => X"137bfbbf",
		16#2cdb# => X"93060000",
		16#2cdc# => X"a30d0102",
		16#2cdd# => X"1306f0ff",
		16#2cde# => X"6308c940",
		16#2cdf# => X"13060b00",
		16#2ce0# => X"b3e59801",
		16#2ce1# => X"137bfbf7",
		16#2ce2# => X"63900540",
		16#2ce3# => X"63080956",
		16#2ce4# => X"13061000",
		16#2ce5# => X"639ec63e",
		16#2ce6# => X"6ff0dfef",
		16#2ce7# => X"93760b01",
		16#2ce8# => X"130c4d00",
		16#2ce9# => X"63860600",
		16#2cea# => X"83280d00",
		16#2ceb# => X"6f000001",
		16#2cec# => X"93760b04",
		16#2ced# => X"63880600",
		16#2cee# => X"83580d00",
		16#2cef# => X"930c0000",
		16#2cf0# => X"6ff09ffa",
		16#2cf1# => X"93760b20",
		16#2cf2# => X"e38006fe",
		16#2cf3# => X"83480d00",
		16#2cf4# => X"6ff0dffe",
		16#2cf5# => X"b786ffff",
		16#2cf6# => X"93c60683",
		16#2cf7# => X"231ed102",
		16#2cf8# => X"83280d00",
		16#2cf9# => X"b7460110",
		16#2cfa# => X"93874690",
		16#2cfb# => X"130c4d00",
		16#2cfc# => X"930c0000",
		16#2cfd# => X"136b2b00",
		16#2cfe# => X"2324f100",
		16#2cff# => X"93062000",
		16#2d00# => X"6ff01ff7",
		16#2d01# => X"a30d0102",
		16#2d02# => X"9306f0ff",
		16#2d03# => X"130c4d00",
		16#2d04# => X"83240d00",
		16#2d05# => X"6308d92a",
		16#2d06# => X"13060900",
		16#2d07# => X"93050000",
		16#2d08# => X"13850400",
		16#2d09# => X"efb09ff5",
		16#2d0a# => X"930c0000",
		16#2d0b# => X"63040500",
		16#2d0c# => X"33099540",
		16#2d0d# => X"138d0c00",
		16#2d0e# => X"63d42c01",
		16#2d0f# => X"130d0900",
		16#2d10# => X"8346b103",
		16#2d11# => X"63840600",
		16#2d12# => X"130d1d00",
		16#2d13# => X"937d2b00",
		16#2d14# => X"63840d00",
		16#2d15# => X"130d2d00",
		16#2d16# => X"93774b08",
		16#2d17# => X"232cf100",
		16#2d18# => X"63940706",
		16#2d19# => X"b386aa41",
		16#2d1a# => X"6350d006",
		16#2d1b# => X"b7470110",
		16#2d1c# => X"93080001",
		16#2d1d# => X"13888735",
		16#2d1e# => X"13037000",
		16#2d1f# => X"03264104",
		16#2d20# => X"23a00b01",
		16#2d21# => X"83258104",
		16#2d22# => X"13061600",
		16#2d23# => X"13858b00",
		16#2d24# => X"63ced848",
		16#2d25# => X"23a2db00",
		16#2d26# => X"b386b600",
		16#2d27# => X"2324d104",
		16#2d28# => X"2322c104",
		16#2d29# => X"93067000",
		16#2d2a# => X"930b0500",
		16#2d2b# => X"63dec600",
		16#2d2c# => X"13060104",
		16#2d2d# => X"93050400",
		16#2d2e# => X"13850900",
		16#2d2f# => X"eff0df89",
		16#2d30# => X"6312055a",
		16#2d31# => X"930bc104",
		16#2d32# => X"8346b103",
		16#2d33# => X"63880604",
		16#2d34# => X"1306b103",
		16#2d35# => X"23a0cb00",
		16#2d36# => X"13061000",
		16#2d37# => X"83264104",
		16#2d38# => X"23a2cb00",
		16#2d39# => X"03268104",
		16#2d3a# => X"93861600",
		16#2d3b# => X"2322d104",
		16#2d3c# => X"13061600",
		16#2d3d# => X"2324c104",
		16#2d3e# => X"13067000",
		16#2d3f# => X"938b8b00",
		16#2d40# => X"635ed600",
		16#2d41# => X"13060104",
		16#2d42# => X"93050400",
		16#2d43# => X"13850900",
		16#2d44# => X"eff09f84",
		16#2d45# => X"63180554",
		16#2d46# => X"930bc104",
		16#2d47# => X"63880d04",
		16#2d48# => X"1306c103",
		16#2d49# => X"23a0cb00",
		16#2d4a# => X"13062000",
		16#2d4b# => X"83264104",
		16#2d4c# => X"23a2cb00",
		16#2d4d# => X"03268104",
		16#2d4e# => X"93861600",
		16#2d4f# => X"2322d104",
		16#2d50# => X"13062600",
		16#2d51# => X"2324c104",
		16#2d52# => X"13067000",
		16#2d53# => X"938b8b00",
		16#2d54# => X"635ed600",
		16#2d55# => X"13060104",
		16#2d56# => X"93050400",
		16#2d57# => X"13850900",
		16#2d58# => X"eff08fff",
		16#2d59# => X"63100550",
		16#2d5a# => X"930bc104",
		16#2d5b# => X"83278101",
		16#2d5c# => X"93060008",
		16#2d5d# => X"6392d706",
		16#2d5e# => X"b38daa41",
		16#2d5f# => X"635eb005",
		16#2d60# => X"13080001",
		16#2d61# => X"93087000",
		16#2d62# => X"83270101",
		16#2d63# => X"83264104",
		16#2d64# => X"03268104",
		16#2d65# => X"23a0fb00",
		16#2d66# => X"93861600",
		16#2d67# => X"93858b00",
		16#2d68# => X"6342b83f",
		16#2d69# => X"23a2bb01",
		16#2d6a# => X"b38dcd00",
		16#2d6b# => X"2324b105",
		16#2d6c# => X"2322d104",
		16#2d6d# => X"13067000",
		16#2d6e# => X"938b0500",
		16#2d6f# => X"635ed600",
		16#2d70# => X"13060104",
		16#2d71# => X"93050400",
		16#2d72# => X"13850900",
		16#2d73# => X"eff0cff8",
		16#2d74# => X"631a0548",
		16#2d75# => X"930bc104",
		16#2d76# => X"b38c2c41",
		16#2d77# => X"635e9005",
		16#2d78# => X"930d0001",
		16#2d79# => X"13087000",
		16#2d7a# => X"83270101",
		16#2d7b# => X"83264104",
		16#2d7c# => X"03268104",
		16#2d7d# => X"23a0fb00",
		16#2d7e# => X"93861600",
		16#2d7f# => X"93858b00",
		16#2d80# => X"63c69d3d",
		16#2d81# => X"23a29b01",
		16#2d82# => X"b38ccc00",
		16#2d83# => X"23249105",
		16#2d84# => X"2322d104",
		16#2d85# => X"13067000",
		16#2d86# => X"938b0500",
		16#2d87# => X"635ed600",
		16#2d88# => X"13060104",
		16#2d89# => X"93050400",
		16#2d8a# => X"13850900",
		16#2d8b# => X"eff0cff2",
		16#2d8c# => X"631a0542",
		16#2d8d# => X"930bc104",
		16#2d8e# => X"83268104",
		16#2d8f# => X"23a22b01",
		16#2d90# => X"23a09b00",
		16#2d91# => X"33892601",
		16#2d92# => X"83264104",
		16#2d93# => X"23242105",
		16#2d94# => X"13067000",
		16#2d95# => X"93861600",
		16#2d96# => X"2322d104",
		16#2d97# => X"13878b00",
		16#2d98# => X"635ed600",
		16#2d99# => X"13060104",
		16#2d9a# => X"93050400",
		16#2d9b# => X"13850900",
		16#2d9c# => X"eff08fee",
		16#2d9d# => X"6318053e",
		16#2d9e# => X"1307c104",
		16#2d9f# => X"93774b00",
		16#2da0# => X"63960738",
		16#2da1# => X"63d4aa01",
		16#2da2# => X"930a0d00",
		16#2da3# => X"83270100",
		16#2da4# => X"b3875701",
		16#2da5# => X"2320f100",
		16#2da6# => X"83278104",
		16#2da7# => X"638c0700",
		16#2da8# => X"13060104",
		16#2da9# => X"93050400",
		16#2daa# => X"13850900",
		16#2dab# => X"eff0cfea",
		16#2dac# => X"631a053a",
		16#2dad# => X"23220104",
		16#2dae# => X"130d0c00",
		16#2daf# => X"930bc104",
		16#2db0# => X"6ff0df8f",
		16#2db1# => X"13850400",
		16#2db2# => X"ef60cf94",
		16#2db3# => X"13090500",
		16#2db4# => X"930c0000",
		16#2db5# => X"6ff01fd6",
		16#2db6# => X"136b0b01",
		16#2db7# => X"93760b02",
		16#2db8# => X"63800602",
		16#2db9# => X"130d7d00",
		16#2dba# => X"137d8dff",
		16#2dbb# => X"83280d00",
		16#2dbc# => X"832c4d00",
		16#2dbd# => X"130c8d00",
		16#2dbe# => X"93061000",
		16#2dbf# => X"6ff05fc7",
		16#2dc0# => X"93760b01",
		16#2dc1# => X"130c4d00",
		16#2dc2# => X"63860600",
		16#2dc3# => X"83280d00",
		16#2dc4# => X"6f000001",
		16#2dc5# => X"93760b04",
		16#2dc6# => X"63880600",
		16#2dc7# => X"83580d00",
		16#2dc8# => X"930c0000",
		16#2dc9# => X"6ff05ffd",
		16#2dca# => X"93760b20",
		16#2dcb# => X"e38006fe",
		16#2dcc# => X"83480d00",
		16#2dcd# => X"6ff0dffe",
		16#2dce# => X"b7460110",
		16#2dcf# => X"93874690",
		16#2dd0# => X"6ff01f94",
		16#2dd1# => X"93760b01",
		16#2dd2# => X"130c4d00",
		16#2dd3# => X"63860600",
		16#2dd4# => X"83280d00",
		16#2dd5# => X"6f000001",
		16#2dd6# => X"93760b04",
		16#2dd7# => X"63880600",
		16#2dd8# => X"83580d00",
		16#2dd9# => X"930c0000",
		16#2dda# => X"6ff09f93",
		16#2ddb# => X"93760b20",
		16#2ddc# => X"e38006fe",
		16#2ddd# => X"83480d00",
		16#2dde# => X"6ff0dffe",
		16#2ddf# => X"13060b00",
		16#2de0# => X"93061000",
		16#2de1# => X"6ff0dfbf",
		16#2de2# => X"13061000",
		16#2de3# => X"e38ec6ae",
		16#2de4# => X"13062000",
		16#2de5# => X"6388c612",
		16#2de6# => X"9306010f",
		16#2de7# => X"9395dc01",
		16#2de8# => X"13f67800",
		16#2de9# => X"93d83800",
		16#2dea# => X"13060603",
		16#2deb# => X"b3e81501",
		16#2dec# => X"93dc3c00",
		16#2ded# => X"a38fc6fe",
		16#2dee# => X"b3e59801",
		16#2def# => X"9384f6ff",
		16#2df0# => X"63960502",
		16#2df1# => X"93751b00",
		16#2df2# => X"638a0500",
		16#2df3# => X"93050003",
		16#2df4# => X"6306b600",
		16#2df5# => X"a38fb4fe",
		16#2df6# => X"9384e6ff",
		16#2df7# => X"9307010f",
		16#2df8# => X"930c0900",
		16#2df9# => X"33899740",
		16#2dfa# => X"6ff0dfc4",
		16#2dfb# => X"93860400",
		16#2dfc# => X"6ff0dffa",
		16#2dfd# => X"93770b40",
		16#2dfe# => X"130d0000",
		16#2dff# => X"130e010f",
		16#2e00# => X"232cf100",
		16#2e01# => X"930d9000",
		16#2e02# => X"13850800",
		16#2e03# => X"1306a000",
		16#2e04# => X"93060000",
		16#2e05# => X"93850c00",
		16#2e06# => X"9304feff",
		16#2e07# => X"2322c103",
		16#2e08# => X"23201103",
		16#2e09# => X"ef20c049",
		16#2e0a# => X"032e4102",
		16#2e0b# => X"83278101",
		16#2e0c# => X"13050503",
		16#2e0d# => X"a30faefe",
		16#2e0e# => X"130d1d00",
		16#2e0f# => X"83280102",
		16#2e10# => X"638c0704",
		16#2e11# => X"83274100",
		16#2e12# => X"83c60700",
		16#2e13# => X"6396a605",
		16#2e14# => X"9307f00f",
		16#2e15# => X"6302fd04",
		16#2e16# => X"63940c00",
		16#2e17# => X"63fe1d03",
		16#2e18# => X"8327c100",
		16#2e19# => X"83254101",
		16#2e1a# => X"23201103",
		16#2e1b# => X"b384f440",
		16#2e1c# => X"13860700",
		16#2e1d# => X"13850400",
		16#2e1e# => X"efd08fd3",
		16#2e1f# => X"83274100",
		16#2e20# => X"130d0000",
		16#2e21# => X"83280102",
		16#2e22# => X"83c61700",
		16#2e23# => X"63860600",
		16#2e24# => X"93871700",
		16#2e25# => X"2322f100",
		16#2e26# => X"13850800",
		16#2e27# => X"93850c00",
		16#2e28# => X"1306a000",
		16#2e29# => X"93060000",
		16#2e2a# => X"ef10d063",
		16#2e2b# => X"938c0500",
		16#2e2c# => X"b3e5a500",
		16#2e2d# => X"93080500",
		16#2e2e# => X"e38205f2",
		16#2e2f# => X"138e0400",
		16#2e30# => X"6ff09ff4",
		16#2e31# => X"9304010f",
		16#2e32# => X"83278100",
		16#2e33# => X"93f6f800",
		16#2e34# => X"9384f4ff",
		16#2e35# => X"b386d700",
		16#2e36# => X"83c60600",
		16#2e37# => X"93d84800",
		16#2e38# => X"2380d400",
		16#2e39# => X"9396cc01",
		16#2e3a# => X"b3e81601",
		16#2e3b# => X"93dc4c00",
		16#2e3c# => X"b3e69801",
		16#2e3d# => X"e39a06fc",
		16#2e3e# => X"6ff05fee",
		16#2e3f# => X"9304010f",
		16#2e40# => X"e39e06ec",
		16#2e41# => X"13761600",
		16#2e42# => X"e30a06ec",
		16#2e43# => X"93060003",
		16#2e44# => X"a307d10e",
		16#2e45# => X"6ff09f98",
		16#2e46# => X"638a0d18",
		16#2e47# => X"2306b109",
		16#2e48# => X"a30d0102",
		16#2e49# => X"130c0d00",
		16#2e4a# => X"6ff0df90",
		16#2e4b# => X"93850501",
		16#2e4c# => X"23a21b01",
		16#2e4d# => X"2324b104",
		16#2e4e# => X"2322c104",
		16#2e4f# => X"635ec302",
		16#2e50# => X"13060104",
		16#2e51# => X"93050400",
		16#2e52# => X"13850900",
		16#2e53# => X"23266102",
		16#2e54# => X"23240103",
		16#2e55# => X"23221103",
		16#2e56# => X"2320d102",
		16#2e57# => X"eff0cfbf",
		16#2e58# => X"63120510",
		16#2e59# => X"0323c102",
		16#2e5a# => X"03288102",
		16#2e5b# => X"83284102",
		16#2e5c# => X"83260102",
		16#2e5d# => X"1305c104",
		16#2e5e# => X"938606ff",
		16#2e5f# => X"930b0500",
		16#2e60# => X"6ff0dfaf",
		16#2e61# => X"13060601",
		16#2e62# => X"23a20b01",
		16#2e63# => X"2324c104",
		16#2e64# => X"2322d104",
		16#2e65# => X"63d6d802",
		16#2e66# => X"13060104",
		16#2e67# => X"93050400",
		16#2e68# => X"13850900",
		16#2e69# => X"23201103",
		16#2e6a# => X"232c0101",
		16#2e6b# => X"eff0cfba",
		16#2e6c# => X"631a050a",
		16#2e6d# => X"83280102",
		16#2e6e# => X"03288101",
		16#2e6f# => X"9305c104",
		16#2e70# => X"938d0dff",
		16#2e71# => X"938b0500",
		16#2e72# => X"6ff01fbc",
		16#2e73# => X"13060601",
		16#2e74# => X"23a2bb01",
		16#2e75# => X"2324c104",
		16#2e76# => X"2322d104",
		16#2e77# => X"6352d802",
		16#2e78# => X"13060104",
		16#2e79# => X"93050400",
		16#2e7a# => X"13850900",
		16#2e7b# => X"232c0101",
		16#2e7c# => X"eff08fb6",
		16#2e7d# => X"63180506",
		16#2e7e# => X"03288101",
		16#2e7f# => X"9305c104",
		16#2e80# => X"938c0cff",
		16#2e81# => X"938b0500",
		16#2e82# => X"6ff01fbe",
		16#2e83# => X"b384aa41",
		16#2e84# => X"e35a90c6",
		16#2e85# => X"b7470110",
		16#2e86# => X"930c0001",
		16#2e87# => X"13898735",
		16#2e88# => X"930d7000",
		16#2e89# => X"83274104",
		16#2e8a# => X"23202701",
		16#2e8b# => X"83268104",
		16#2e8c# => X"93871700",
		16#2e8d# => X"63c09c04",
		16#2e8e# => X"23229700",
		16#2e8f# => X"b384d400",
		16#2e90# => X"23249104",
		16#2e91# => X"2322f104",
		16#2e92# => X"13077000",
		16#2e93# => X"e35cf7c2",
		16#2e94# => X"13060104",
		16#2e95# => X"93050400",
		16#2e96# => X"13850900",
		16#2e97# => X"eff0cfaf",
		16#2e98# => X"e30205c2",
		16#2e99# => X"8357c400",
		16#2e9a# => X"93f70704",
		16#2e9b# => X"638a07ca",
		16#2e9c# => X"6ff00fd0",
		16#2e9d# => X"93860601",
		16#2e9e# => X"23229701",
		16#2e9f# => X"2324d104",
		16#2ea0# => X"2322f104",
		16#2ea1# => X"13078700",
		16#2ea2# => X"63defd00",
		16#2ea3# => X"13060104",
		16#2ea4# => X"93050400",
		16#2ea5# => X"13850900",
		16#2ea6# => X"eff00fac",
		16#2ea7# => X"e31405fc",
		16#2ea8# => X"1307c104",
		16#2ea9# => X"938404ff",
		16#2eaa# => X"6ff0dff7",
		16#2eab# => X"83278104",
		16#2eac# => X"e38a07fa",
		16#2ead# => X"13060104",
		16#2eae# => X"93050400",
		16#2eaf# => X"13850900",
		16#2eb0# => X"eff08fa9",
		16#2eb1# => X"6ff01ffa",
		16#2eb2# => X"93060600",
		16#2eb3# => X"13860500",
		16#2eb4# => X"93050500",
		16#2eb5# => X"03a5c181",
		16#2eb6# => X"6ff00fb8",
		16#2eb7# => X"83d7c500",
		16#2eb8# => X"130101b8",
		16#2eb9# => X"232c8146",
		16#2eba# => X"93f7d7ff",
		16#2ebb# => X"231af100",
		16#2ebc# => X"83a74506",
		16#2ebd# => X"13840500",
		16#2ebe# => X"232a9146",
		16#2ebf# => X"2326f106",
		16#2ec0# => X"83d7e500",
		16#2ec1# => X"23282147",
		16#2ec2# => X"232e1146",
		16#2ec3# => X"231bf100",
		16#2ec4# => X"83a7c501",
		16#2ec5# => X"13090500",
		16#2ec6# => X"23200102",
		16#2ec7# => X"2322f102",
		16#2ec8# => X"83a74502",
		16#2ec9# => X"93058100",
		16#2eca# => X"2326f102",
		16#2ecb# => X"93070107",
		16#2ecc# => X"2324f100",
		16#2ecd# => X"232cf100",
		16#2ece# => X"93070040",
		16#2ecf# => X"2328f100",
		16#2ed0# => X"232ef100",
		16#2ed1# => X"eff04fb1",
		16#2ed2# => X"93040500",
		16#2ed3# => X"634c0500",
		16#2ed4# => X"93058100",
		16#2ed5# => X"13050900",
		16#2ed6# => X"ef804f9f",
		16#2ed7# => X"63040500",
		16#2ed8# => X"9304f0ff",
		16#2ed9# => X"83574101",
		16#2eda# => X"93f70704",
		16#2edb# => X"63880700",
		16#2edc# => X"8357c400",
		16#2edd# => X"93e70704",
		16#2ede# => X"2316f400",
		16#2edf# => X"8320c147",
		16#2ee0# => X"03248147",
		16#2ee1# => X"13850400",
		16#2ee2# => X"03290147",
		16#2ee3# => X"83244147",
		16#2ee4# => X"13010148",
		16#2ee5# => X"67800000",
		16#2ee6# => X"83a7c181",
		16#2ee7# => X"83a74703",
		16#2ee8# => X"63960700",
		16#2ee9# => X"b7570110",
		16#2eea# => X"938707ca",
		16#2eeb# => X"03a3070e",
		16#2eec# => X"67000300",
		16#2eed# => X"63840502",
		16#2eee# => X"9307f00f",
		16#2eef# => X"63fac700",
		16#2ef0# => X"9307a008",
		16#2ef1# => X"2320f500",
		16#2ef2# => X"1305f0ff",
		16#2ef3# => X"67800000",
		16#2ef4# => X"2380c500",
		16#2ef5# => X"13051000",
		16#2ef6# => X"67800000",
		16#2ef7# => X"13050000",
		16#2ef8# => X"67800000",
		16#2ef9# => X"130101ff",
		16#2efa# => X"23248100",
		16#2efb# => X"23229100",
		16#2efc# => X"37840110",
		16#2efd# => X"93040500",
		16#2efe# => X"13850500",
		16#2eff# => X"93050600",
		16#2f00# => X"13860600",
		16#2f01# => X"23261100",
		16#2f02# => X"232204aa",
		16#2f03# => X"ef10900e",
		16#2f04# => X"9307f0ff",
		16#2f05# => X"6318f500",
		16#2f06# => X"832744aa",
		16#2f07# => X"63840700",
		16#2f08# => X"23a0f400",
		16#2f09# => X"8320c100",
		16#2f0a# => X"03248100",
		16#2f0b# => X"83244100",
		16#2f0c# => X"13010101",
		16#2f0d# => X"67800000",
		16#2f0e# => X"130101ff",
		16#2f0f# => X"23248100",
		16#2f10# => X"13040500",
		16#2f11# => X"13850500",
		16#2f12# => X"93050600",
		16#2f13# => X"23261100",
		16#2f14# => X"ef60101e",
		16#2f15# => X"93050500",
		16#2f16# => X"13050400",
		16#2f17# => X"efb0cf85",
		16#2f18# => X"13040500",
		16#2f19# => X"63020504",
		16#2f1a# => X"0326c5ff",
		16#2f1b# => X"13074002",
		16#2f1c# => X"1376c6ff",
		16#2f1d# => X"1306c6ff",
		16#2f1e# => X"6362c706",
		16#2f1f# => X"93063001",
		16#2f20# => X"93070500",
		16#2f21# => X"63fcc600",
		16#2f22# => X"23200500",
		16#2f23# => X"23220500",
		16#2f24# => X"9307b001",
		16#2f25# => X"63e4c702",
		16#2f26# => X"93078500",
		16#2f27# => X"23a00700",
		16#2f28# => X"23a20700",
		16#2f29# => X"23a40700",
		16#2f2a# => X"13050400",
		16#2f2b# => X"8320c100",
		16#2f2c# => X"03248100",
		16#2f2d# => X"13010101",
		16#2f2e# => X"67800000",
		16#2f2f# => X"23240500",
		16#2f30# => X"23260500",
		16#2f31# => X"93070501",
		16#2f32# => X"e31ae6fc",
		16#2f33# => X"23280500",
		16#2f34# => X"93078501",
		16#2f35# => X"232a0500",
		16#2f36# => X"6ff05ffc",
		16#2f37# => X"93050000",
		16#2f38# => X"efb0cfff",
		16#2f39# => X"6ff05ffc",
		16#2f3a# => X"130101ff",
		16#2f3b# => X"23248100",
		16#2f3c# => X"23229100",
		16#2f3d# => X"37840110",
		16#2f3e# => X"93040500",
		16#2f3f# => X"13850500",
		16#2f40# => X"23261100",
		16#2f41# => X"232204aa",
		16#2f42# => X"ef109006",
		16#2f43# => X"9307f0ff",
		16#2f44# => X"6318f500",
		16#2f45# => X"832744aa",
		16#2f46# => X"63840700",
		16#2f47# => X"23a0f400",
		16#2f48# => X"8320c100",
		16#2f49# => X"03248100",
		16#2f4a# => X"83244100",
		16#2f4b# => X"13010101",
		16#2f4c# => X"67800000",
		16#2f4d# => X"130101ff",
		16#2f4e# => X"23261100",
		16#2f4f# => X"23248100",
		16#2f50# => X"23229100",
		16#2f51# => X"23202101",
		16#2f52# => X"63920502",
		16#2f53# => X"13090000",
		16#2f54# => X"8320c100",
		16#2f55# => X"03248100",
		16#2f56# => X"13050900",
		16#2f57# => X"83244100",
		16#2f58# => X"03290100",
		16#2f59# => X"13010101",
		16#2f5a# => X"67800000",
		16#2f5b# => X"93040500",
		16#2f5c# => X"13840500",
		16#2f5d# => X"63080500",
		16#2f5e# => X"83278503",
		16#2f5f# => X"63940700",
		16#2f60# => X"ef808f96",
		16#2f61# => X"8317c400",
		16#2f62# => X"e38207fc",
		16#2f63# => X"93050400",
		16#2f64# => X"13850400",
		16#2f65# => X"ef701fdb",
		16#2f66# => X"8327c402",
		16#2f67# => X"13090500",
		16#2f68# => X"638c0700",
		16#2f69# => X"8325c401",
		16#2f6a# => X"13850400",
		16#2f6b# => X"e7800700",
		16#2f6c# => X"63540500",
		16#2f6d# => X"1309f0ff",
		16#2f6e# => X"8357c400",
		16#2f6f# => X"93f70708",
		16#2f70# => X"63880700",
		16#2f71# => X"83250401",
		16#2f72# => X"13850400",
		16#2f73# => X"ef800fbd",
		16#2f74# => X"83250403",
		16#2f75# => X"638c0500",
		16#2f76# => X"93070404",
		16#2f77# => X"6386f500",
		16#2f78# => X"13850400",
		16#2f79# => X"ef808fbb",
		16#2f7a# => X"23280402",
		16#2f7b# => X"83254404",
		16#2f7c# => X"63880500",
		16#2f7d# => X"13850400",
		16#2f7e# => X"ef804fba",
		16#2f7f# => X"23220404",
		16#2f80# => X"ef804fa5",
		16#2f81# => X"23160400",
		16#2f82# => X"ef800fa5",
		16#2f83# => X"6ff05ff4",
		16#2f84# => X"93050500",
		16#2f85# => X"03a5c181",
		16#2f86# => X"6ff0dff1",
		16#2f87# => X"130101fd",
		16#2f88# => X"23248102",
		16#2f89# => X"23229102",
		16#2f8a# => X"232c4101",
		16#2f8b# => X"23261102",
		16#2f8c# => X"23202103",
		16#2f8d# => X"232e3101",
		16#2f8e# => X"232a5101",
		16#2f8f# => X"23286101",
		16#2f90# => X"130a0500",
		16#2f91# => X"93840500",
		16#2f92# => X"13040600",
		16#2f93# => X"efa01fc9",
		16#2f94# => X"93071000",
		16#2f95# => X"631af504",
		16#2f96# => X"9387f4ff",
		16#2f97# => X"1307e00f",
		16#2f98# => X"6364f704",
		16#2f99# => X"23069100",
		16#2f9a# => X"93091000",
		16#2f9b# => X"13090000",
		16#2f9c# => X"930af0ff",
		16#2f9d# => X"130ba000",
		16#2f9e# => X"63123907",
		16#2f9f# => X"13850400",
		16#2fa0# => X"8320c102",
		16#2fa1# => X"03248102",
		16#2fa2# => X"83244102",
		16#2fa3# => X"03290102",
		16#2fa4# => X"8329c101",
		16#2fa5# => X"032a8101",
		16#2fa6# => X"832a4101",
		16#2fa7# => X"032b0101",
		16#2fa8# => X"13010103",
		16#2fa9# => X"67800000",
		16#2faa# => X"9306c405",
		16#2fab# => X"13860400",
		16#2fac# => X"9305c100",
		16#2fad# => X"13050a00",
		16#2fae# => X"ef104016",
		16#2faf# => X"9307f0ff",
		16#2fb0# => X"93090500",
		16#2fb1# => X"e314f5fa",
		16#2fb2# => X"8357c400",
		16#2fb3# => X"93e70704",
		16#2fb4# => X"2316f400",
		16#2fb5# => X"1305f0ff",
		16#2fb6# => X"6ff09ffa",
		16#2fb7# => X"9307c100",
		16#2fb8# => X"b3872701",
		16#2fb9# => X"83c50700",
		16#2fba# => X"83278400",
		16#2fbb# => X"9387f7ff",
		16#2fbc# => X"2324f400",
		16#2fbd# => X"63d80700",
		16#2fbe# => X"03278401",
		16#2fbf# => X"63c0e702",
		16#2fc0# => X"638e6501",
		16#2fc1# => X"83270400",
		16#2fc2# => X"13871700",
		16#2fc3# => X"2320e400",
		16#2fc4# => X"2380b700",
		16#2fc5# => X"13091900",
		16#2fc6# => X"6ff01ff6",
		16#2fc7# => X"13060400",
		16#2fc8# => X"13050a00",
		16#2fc9# => X"ef70df9a",
		16#2fca# => X"e31655ff",
		16#2fcb# => X"6ff09ffa",
		16#2fcc# => X"8317c600",
		16#2fcd# => X"13972701",
		16#2fce# => X"63400702",
		16#2fcf# => X"03274606",
		16#2fd0# => X"b7260000",
		16#2fd1# => X"b3e7d700",
		16#2fd2# => X"2316f600",
		16#2fd3# => X"b7270000",
		16#2fd4# => X"b367f700",
		16#2fd5# => X"2322f606",
		16#2fd6# => X"6ff05fec",
		16#2fd7# => X"130101fe",
		16#2fd8# => X"232c8100",
		16#2fd9# => X"03a4c181",
		16#2fda# => X"232a9100",
		16#2fdb# => X"232e1100",
		16#2fdc# => X"93040500",
		16#2fdd# => X"13860500",
		16#2fde# => X"630e0400",
		16#2fdf# => X"83278403",
		16#2fe0# => X"639a0700",
		16#2fe1# => X"13050400",
		16#2fe2# => X"2326b100",
		16#2fe3# => X"ef70dff5",
		16#2fe4# => X"0326c100",
		16#2fe5# => X"13050400",
		16#2fe6# => X"03248101",
		16#2fe7# => X"8320c101",
		16#2fe8# => X"93850400",
		16#2fe9# => X"83244101",
		16#2fea# => X"13010102",
		16#2feb# => X"6ff05ff8",
		16#2fec# => X"130101ff",
		16#2fed# => X"23248100",
		16#2fee# => X"23229100",
		16#2fef# => X"37840110",
		16#2ff0# => X"93040500",
		16#2ff1# => X"13850500",
		16#2ff2# => X"93050600",
		16#2ff3# => X"23261100",
		16#2ff4# => X"232204aa",
		16#2ff5# => X"ef10405a",
		16#2ff6# => X"9307f0ff",
		16#2ff7# => X"6318f500",
		16#2ff8# => X"832744aa",
		16#2ff9# => X"63840700",
		16#2ffa# => X"23a0f400",
		16#2ffb# => X"8320c100",
		16#2ffc# => X"03248100",
		16#2ffd# => X"83244100",
		16#2ffe# => X"13010101",
		16#2fff# => X"67800000",
		16#3000# => X"130101ff",
		16#3001# => X"23248100",
		16#3002# => X"23229100",
		16#3003# => X"37840110",
		16#3004# => X"93040500",
		16#3005# => X"13850500",
		16#3006# => X"23261100",
		16#3007# => X"232204aa",
		16#3008# => X"ef108056",
		16#3009# => X"9307f0ff",
		16#300a# => X"6318f500",
		16#300b# => X"832744aa",
		16#300c# => X"63840700",
		16#300d# => X"23a0f400",
		16#300e# => X"8320c100",
		16#300f# => X"03248100",
		16#3010# => X"83244100",
		16#3011# => X"13010101",
		16#3012# => X"67800000",
		16#3013# => X"130101ff",
		16#3014# => X"23248100",
		16#3015# => X"23229100",
		16#3016# => X"37840110",
		16#3017# => X"93040500",
		16#3018# => X"13850500",
		16#3019# => X"93050600",
		16#301a# => X"13860600",
		16#301b# => X"23261100",
		16#301c# => X"232204aa",
		16#301d# => X"ef10c051",
		16#301e# => X"9307f0ff",
		16#301f# => X"6318f500",
		16#3020# => X"832744aa",
		16#3021# => X"63840700",
		16#3022# => X"23a0f400",
		16#3023# => X"8320c100",
		16#3024# => X"03248100",
		16#3025# => X"83244100",
		16#3026# => X"13010101",
		16#3027# => X"67800000",
		16#3028# => X"130101ff",
		16#3029# => X"23248100",
		16#302a# => X"23229100",
		16#302b# => X"37840110",
		16#302c# => X"93040500",
		16#302d# => X"13850500",
		16#302e# => X"93050600",
		16#302f# => X"13860600",
		16#3030# => X"23261100",
		16#3031# => X"232204aa",
		16#3032# => X"ef10403d",
		16#3033# => X"9307f0ff",
		16#3034# => X"6318f500",
		16#3035# => X"832744aa",
		16#3036# => X"63840700",
		16#3037# => X"23a0f400",
		16#3038# => X"8320c100",
		16#3039# => X"03248100",
		16#303a# => X"83244100",
		16#303b# => X"13010101",
		16#303c# => X"67800000",
		16#303d# => X"130101ff",
		16#303e# => X"23248100",
		16#303f# => X"13840500",
		16#3040# => X"83a50500",
		16#3041# => X"23229100",
		16#3042# => X"23261100",
		16#3043# => X"93040500",
		16#3044# => X"63840500",
		16#3045# => X"eff01ffe",
		16#3046# => X"93050400",
		16#3047# => X"03248100",
		16#3048# => X"8320c100",
		16#3049# => X"13850400",
		16#304a# => X"83244100",
		16#304b# => X"13010101",
		16#304c# => X"6f80cf86",
		16#304d# => X"83a7c181",
		16#304e# => X"6382a710",
		16#304f# => X"8327c504",
		16#3050# => X"130101fe",
		16#3051# => X"232c8100",
		16#3052# => X"232a9100",
		16#3053# => X"23282101",
		16#3054# => X"232e1100",
		16#3055# => X"23263101",
		16#3056# => X"13040500",
		16#3057# => X"93040000",
		16#3058# => X"13090008",
		16#3059# => X"63940704",
		16#305a# => X"83250404",
		16#305b# => X"63860500",
		16#305c# => X"13050400",
		16#305d# => X"ef808f82",
		16#305e# => X"83258414",
		16#305f# => X"638c0504",
		16#3060# => X"9304c414",
		16#3061# => X"63889504",
		16#3062# => X"03a90500",
		16#3063# => X"13050400",
		16#3064# => X"ef80cf80",
		16#3065# => X"93050900",
		16#3066# => X"6ff0dffe",
		16#3067# => X"b3859500",
		16#3068# => X"83a50500",
		16#3069# => X"639e0500",
		16#306a# => X"93844400",
		16#306b# => X"8325c404",
		16#306c# => X"e39624ff",
		16#306d# => X"13050400",
		16#306e# => X"ef705ffe",
		16#306f# => X"6ff0dffa",
		16#3070# => X"83a90500",
		16#3071# => X"13050400",
		16#3072# => X"ef705ffd",
		16#3073# => X"93850900",
		16#3074# => X"6ff05ffd",
		16#3075# => X"83254405",
		16#3076# => X"63860500",
		16#3077# => X"13050400",
		16#3078# => X"ef70dffb",
		16#3079# => X"83278403",
		16#307a# => X"638c0702",
		16#307b# => X"8327c403",
		16#307c# => X"13050400",
		16#307d# => X"e7800700",
		16#307e# => X"8325042e",
		16#307f# => X"63820502",
		16#3080# => X"13050400",
		16#3081# => X"03248101",
		16#3082# => X"8320c101",
		16#3083# => X"83244101",
		16#3084# => X"03290101",
		16#3085# => X"8329c100",
		16#3086# => X"13010102",
		16#3087# => X"6ff09fed",
		16#3088# => X"8320c101",
		16#3089# => X"03248101",
		16#308a# => X"83244101",
		16#308b# => X"03290101",
		16#308c# => X"8329c100",
		16#308d# => X"13010102",
		16#308e# => X"67800000",
		16#308f# => X"67800000",
		16#3090# => X"83278600",
		16#3091# => X"130101fd",
		16#3092# => X"232e3101",
		16#3093# => X"23261102",
		16#3094# => X"23248102",
		16#3095# => X"23229102",
		16#3096# => X"23202103",
		16#3097# => X"232c4101",
		16#3098# => X"232a5101",
		16#3099# => X"23286101",
		16#309a# => X"23267101",
		16#309b# => X"23248101",
		16#309c# => X"23229101",
		16#309d# => X"93090600",
		16#309e# => X"63860712",
		16#309f# => X"032b0600",
		16#30a0# => X"930a0500",
		16#30a1# => X"13840500",
		16#30a2# => X"930b0000",
		16#30a3# => X"13090000",
		16#30a4# => X"63060908",
		16#30a5# => X"032a8400",
		16#30a6# => X"6366490d",
		16#30a7# => X"835cc400",
		16#30a8# => X"93f70c48",
		16#30a9# => X"6380070c",
		16#30aa# => X"03254401",
		16#30ab# => X"83240400",
		16#30ac# => X"032a0401",
		16#30ad# => X"93053000",
		16#30ae# => X"ef608037",
		16#30af# => X"338c4441",
		16#30b0# => X"9354f501",
		16#30b1# => X"b384a400",
		16#30b2# => X"93071c00",
		16#30b3# => X"93d41440",
		16#30b4# => X"b3872701",
		16#30b5# => X"63f4f400",
		16#30b6# => X"93840700",
		16#30b7# => X"93fc0c40",
		16#30b8# => X"63800c10",
		16#30b9# => X"93850400",
		16#30ba# => X"13850a00",
		16#30bb# => X"efa0df9c",
		16#30bc# => X"130a0500",
		16#30bd# => X"631c0502",
		16#30be# => X"9307c000",
		16#30bf# => X"23a0fa00",
		16#30c0# => X"8357c400",
		16#30c1# => X"1305f0ff",
		16#30c2# => X"93e70704",
		16#30c3# => X"2316f400",
		16#30c4# => X"23a40900",
		16#30c5# => X"23a20900",
		16#30c6# => X"6f004009",
		16#30c7# => X"832b0b00",
		16#30c8# => X"03294b00",
		16#30c9# => X"130b8b00",
		16#30ca# => X"6ff09ff6",
		16#30cb# => X"83250401",
		16#30cc# => X"13060c00",
		16#30cd# => X"efb0cf86",
		16#30ce# => X"8357c400",
		16#30cf# => X"93f7f7b7",
		16#30d0# => X"93e70708",
		16#30d1# => X"2316f400",
		16#30d2# => X"23284401",
		16#30d3# => X"232a9400",
		16#30d4# => X"330a8a01",
		16#30d5# => X"b3848441",
		16#30d6# => X"23204401",
		16#30d7# => X"23249400",
		16#30d8# => X"130a0900",
		16#30d9# => X"63744901",
		16#30da# => X"130a0900",
		16#30db# => X"03250400",
		16#30dc# => X"13060a00",
		16#30dd# => X"93850b00",
		16#30de# => X"efb00f91",
		16#30df# => X"83278400",
		16#30e0# => X"b3874741",
		16#30e1# => X"2324f400",
		16#30e2# => X"83270400",
		16#30e3# => X"338a4701",
		16#30e4# => X"83a78900",
		16#30e5# => X"23204401",
		16#30e6# => X"33892741",
		16#30e7# => X"23a42901",
		16#30e8# => X"e31e09f6",
		16#30e9# => X"23a20900",
		16#30ea# => X"13050000",
		16#30eb# => X"8320c102",
		16#30ec# => X"03248102",
		16#30ed# => X"83244102",
		16#30ee# => X"03290102",
		16#30ef# => X"8329c101",
		16#30f0# => X"032a8101",
		16#30f1# => X"832a4101",
		16#30f2# => X"032b0101",
		16#30f3# => X"832bc100",
		16#30f4# => X"032c8100",
		16#30f5# => X"832c4100",
		16#30f6# => X"13010103",
		16#30f7# => X"67800000",
		16#30f8# => X"93050a00",
		16#30f9# => X"13860400",
		16#30fa# => X"13850a00",
		16#30fb# => X"efc04f94",
		16#30fc# => X"130a0500",
		16#30fd# => X"e31a05f4",
		16#30fe# => X"83250401",
		16#30ff# => X"13850a00",
		16#3100# => X"ef70dfd9",
		16#3101# => X"6ff05fef",
		16#3102# => X"83d7c500",
		16#3103# => X"130101ed",
		16#3104# => X"23202113",
		16#3105# => X"232e3111",
		16#3106# => X"232c4111",
		16#3107# => X"2320a111",
		16#3108# => X"23261112",
		16#3109# => X"23248112",
		16#310a# => X"23229112",
		16#310b# => X"232a5111",
		16#310c# => X"23286111",
		16#310d# => X"23267111",
		16#310e# => X"23248111",
		16#310f# => X"23229111",
		16#3110# => X"232eb10f",
		16#3111# => X"93f70708",
		16#3112# => X"130a0500",
		16#3113# => X"13890500",
		16#3114# => X"93090600",
		16#3115# => X"138d0600",
		16#3116# => X"638e0702",
		16#3117# => X"83a70501",
		16#3118# => X"639a0702",
		16#3119# => X"93050004",
		16#311a# => X"efa01f85",
		16#311b# => X"2320a900",
		16#311c# => X"2328a900",
		16#311d# => X"631c0500",
		16#311e# => X"9307c000",
		16#311f# => X"2320fa00",
		16#3120# => X"9307f0ff",
		16#3121# => X"2320f100",
		16#3122# => X"6f001030",
		16#3123# => X"93070004",
		16#3124# => X"232af900",
		16#3125# => X"9307c104",
		16#3126# => X"2320f104",
		16#3127# => X"938b0700",
		16#3128# => X"b7470110",
		16#3129# => X"9387c747",
		16#312a# => X"232ef100",
		16#312b# => X"b7470110",
		16#312c# => X"9387875f",
		16#312d# => X"23240104",
		16#312e# => X"23220104",
		16#312f# => X"23240100",
		16#3130# => X"23220100",
		16#3131# => X"23260100",
		16#3132# => X"232a0100",
		16#3133# => X"23200100",
		16#3134# => X"2328f100",
		16#3135# => X"13840900",
		16#3136# => X"93065002",
		16#3137# => X"83470400",
		16#3138# => X"63840700",
		16#3139# => X"6392d70a",
		16#313a# => X"b3043441",
		16#313b# => X"638a0404",
		16#313c# => X"83278104",
		16#313d# => X"23a03b01",
		16#313e# => X"23a29b00",
		16#313f# => X"b3879700",
		16#3140# => X"2324f104",
		16#3141# => X"83274104",
		16#3142# => X"93067000",
		16#3143# => X"938b8b00",
		16#3144# => X"93871700",
		16#3145# => X"2322f104",
		16#3146# => X"63def600",
		16#3147# => X"13060104",
		16#3148# => X"93050900",
		16#3149# => X"13050a00",
		16#314a# => X"eff09fd1",
		16#314b# => X"e3180524",
		16#314c# => X"930bc104",
		16#314d# => X"83270100",
		16#314e# => X"b3879700",
		16#314f# => X"2320f100",
		16#3150# => X"83470400",
		16#3151# => X"e38e072a",
		16#3152# => X"93091400",
		16#3153# => X"a30d0102",
		16#3154# => X"9304f0ff",
		16#3155# => X"930a0000",
		16#3156# => X"130b0000",
		16#3157# => X"13049000",
		16#3158# => X"930ca005",
		16#3159# => X"83cd0900",
		16#315a# => X"93891900",
		16#315b# => X"93860dfe",
		16#315c# => X"e3e0dc0c",
		16#315d# => X"8327c101",
		16#315e# => X"93962600",
		16#315f# => X"b386f600",
		16#3160# => X"83a60600",
		16#3161# => X"67800600",
		16#3162# => X"13041400",
		16#3163# => X"6ff01ff5",
		16#3164# => X"b7460110",
		16#3165# => X"93878691",
		16#3166# => X"2324f100",
		16#3167# => X"93760b02",
		16#3168# => X"638e066a",
		16#3169# => X"130d7d00",
		16#316a# => X"137d8dff",
		16#316b# => X"83280d00",
		16#316c# => X"832c4d00",
		16#316d# => X"130c8d00",
		16#316e# => X"93761b00",
		16#316f# => X"638e0600",
		16#3170# => X"b3e69801",
		16#3171# => X"638a0600",
		16#3172# => X"93060003",
		16#3173# => X"230ed102",
		16#3174# => X"a30eb103",
		16#3175# => X"136b2b00",
		16#3176# => X"137bfbbf",
		16#3177# => X"6f008033",
		16#3178# => X"13050a00",
		16#3179# => X"efa0cfc4",
		16#317a# => X"83274500",
		16#317b# => X"13850700",
		16#317c# => X"232af100",
		16#317d# => X"ef500fa2",
		16#317e# => X"2326a100",
		16#317f# => X"13050a00",
		16#3180# => X"efa00fc3",
		16#3181# => X"83278500",
		16#3182# => X"2322f100",
		16#3183# => X"8327c100",
		16#3184# => X"e38807f4",
		16#3185# => X"83274100",
		16#3186# => X"e38407f4",
		16#3187# => X"83c60700",
		16#3188# => X"e38006f4",
		16#3189# => X"136b0b40",
		16#318a# => X"6ff09ff3",
		16#318b# => X"8346b103",
		16#318c# => X"e39806f2",
		16#318d# => X"93060002",
		16#318e# => X"a30dd102",
		16#318f# => X"6ff05ff2",
		16#3190# => X"136b1b00",
		16#3191# => X"6ff0dff1",
		16#3192# => X"832a0d00",
		16#3193# => X"130d4d00",
		16#3194# => X"e3d80af0",
		16#3195# => X"b30a5041",
		16#3196# => X"136b4b00",
		16#3197# => X"6ff05ff0",
		16#3198# => X"9306b002",
		16#3199# => X"6ff05ffd",
		16#319a# => X"83cd0900",
		16#319b# => X"9307a002",
		16#319c# => X"138c1900",
		16#319d# => X"6394fd04",
		16#319e# => X"83240d00",
		16#319f# => X"13064d00",
		16#31a0# => X"63d40400",
		16#31a1# => X"9304f0ff",
		16#31a2# => X"130d0600",
		16#31a3# => X"93090c00",
		16#31a4# => X"6ff01fed",
		16#31a5# => X"13850400",
		16#31a6# => X"9305a000",
		16#31a7# => X"130c1c00",
		16#31a8# => X"ef501079",
		16#31a9# => X"834dfcff",
		16#31aa# => X"b3043501",
		16#31ab# => X"93890dfd",
		16#31ac# => X"e37234ff",
		16#31ad# => X"93090c00",
		16#31ae# => X"6ff05feb",
		16#31af# => X"93040000",
		16#31b0# => X"6ff0dffe",
		16#31b1# => X"136b0b08",
		16#31b2# => X"6ff09fe9",
		16#31b3# => X"138c0900",
		16#31b4# => X"930a0000",
		16#31b5# => X"13850a00",
		16#31b6# => X"9305a000",
		16#31b7# => X"130c1c00",
		16#31b8# => X"ef501075",
		16#31b9# => X"938a0dfd",
		16#31ba# => X"834dfcff",
		16#31bb# => X"b38aaa00",
		16#31bc# => X"13860dfd",
		16#31bd# => X"e370c4fe",
		16#31be# => X"6ff0dffb",
		16#31bf# => X"03c60900",
		16#31c0# => X"93068006",
		16#31c1# => X"6318d600",
		16#31c2# => X"93891900",
		16#31c3# => X"136b0b20",
		16#31c4# => X"6ff01fe5",
		16#31c5# => X"136b0b04",
		16#31c6# => X"6ff09fe4",
		16#31c7# => X"03c60900",
		16#31c8# => X"9306c006",
		16#31c9# => X"6318d600",
		16#31ca# => X"93891900",
		16#31cb# => X"136b0b02",
		16#31cc# => X"6ff01fe3",
		16#31cd# => X"136b0b01",
		16#31ce# => X"6ff09fe2",
		16#31cf# => X"83260d00",
		16#31d0# => X"130c4d00",
		16#31d1# => X"a30d0102",
		16#31d2# => X"2306d108",
		16#31d3# => X"93041000",
		16#31d4# => X"930c0000",
		16#31d5# => X"1304c108",
		16#31d6# => X"6f00401f",
		16#31d7# => X"136b0b01",
		16#31d8# => X"93760b02",
		16#31d9# => X"638c0604",
		16#31da# => X"130d7d00",
		16#31db# => X"137d8dff",
		16#31dc# => X"83280d00",
		16#31dd# => X"832c4d00",
		16#31de# => X"130c8d00",
		16#31df# => X"63de0c00",
		16#31e0# => X"b3081041",
		16#31e1# => X"b3361001",
		16#31e2# => X"33039041",
		16#31e3# => X"b30cd340",
		16#31e4# => X"9306d002",
		16#31e5# => X"a30dd102",
		16#31e6# => X"9306f0ff",
		16#31e7# => X"639cd44e",
		16#31e8# => X"63960c56",
		16#31e9# => X"93069000",
		16#31ea# => X"63e21657",
		16#31eb# => X"93880803",
		16#31ec# => X"a307110f",
		16#31ed# => X"1304f10e",
		16#31ee# => X"6f00c053",
		16#31ef# => X"93760b01",
		16#31f0# => X"130c4d00",
		16#31f1# => X"63880600",
		16#31f2# => X"83280d00",
		16#31f3# => X"93dcf841",
		16#31f4# => X"6ff0dffa",
		16#31f5# => X"93760b04",
		16#31f6# => X"83280d00",
		16#31f7# => X"63880600",
		16#31f8# => X"93980801",
		16#31f9# => X"93d80841",
		16#31fa# => X"6ff05ffe",
		16#31fb# => X"93760b20",
		16#31fc# => X"e38e06fc",
		16#31fd# => X"93988801",
		16#31fe# => X"93d88841",
		16#31ff# => X"6ff01ffd",
		16#3200# => X"13760b02",
		16#3201# => X"83260d00",
		16#3202# => X"130d4d00",
		16#3203# => X"630c0600",
		16#3204# => X"83270100",
		16#3205# => X"23a0f600",
		16#3206# => X"93d7f741",
		16#3207# => X"23a2f600",
		16#3208# => X"6ff05fcb",
		16#3209# => X"13760b01",
		16#320a# => X"63080600",
		16#320b# => X"83270100",
		16#320c# => X"23a0f600",
		16#320d# => X"6ff01fca",
		16#320e# => X"13760b04",
		16#320f# => X"63080600",
		16#3210# => X"83570100",
		16#3211# => X"2390f600",
		16#3212# => X"6ff0dfc8",
		16#3213# => X"93770b20",
		16#3214# => X"e38e07fc",
		16#3215# => X"83470100",
		16#3216# => X"2380f600",
		16#3217# => X"6ff09fc7",
		16#3218# => X"136b0b01",
		16#3219# => X"93760b02",
		16#321a# => X"63860604",
		16#321b# => X"130d7d00",
		16#321c# => X"137d8dff",
		16#321d# => X"83280d00",
		16#321e# => X"832c4d00",
		16#321f# => X"130c8d00",
		16#3220# => X"137bfbbf",
		16#3221# => X"93060000",
		16#3222# => X"a30d0102",
		16#3223# => X"1306f0ff",
		16#3224# => X"6388c440",
		16#3225# => X"13060b00",
		16#3226# => X"b3e59801",
		16#3227# => X"137bfbf7",
		16#3228# => X"63900540",
		16#3229# => X"63880456",
		16#322a# => X"13061000",
		16#322b# => X"639ec63e",
		16#322c# => X"6ff0dfef",
		16#322d# => X"93760b01",
		16#322e# => X"130c4d00",
		16#322f# => X"63860600",
		16#3230# => X"83280d00",
		16#3231# => X"6f000001",
		16#3232# => X"93760b04",
		16#3233# => X"63880600",
		16#3234# => X"83580d00",
		16#3235# => X"930c0000",
		16#3236# => X"6ff09ffa",
		16#3237# => X"93760b20",
		16#3238# => X"e38006fe",
		16#3239# => X"83480d00",
		16#323a# => X"6ff0dffe",
		16#323b# => X"b786ffff",
		16#323c# => X"93c60683",
		16#323d# => X"231ed102",
		16#323e# => X"83280d00",
		16#323f# => X"b7460110",
		16#3240# => X"93874690",
		16#3241# => X"130c4d00",
		16#3242# => X"930c0000",
		16#3243# => X"136b2b00",
		16#3244# => X"2324f100",
		16#3245# => X"93062000",
		16#3246# => X"6ff01ff7",
		16#3247# => X"a30d0102",
		16#3248# => X"9306f0ff",
		16#3249# => X"130c4d00",
		16#324a# => X"03240d00",
		16#324b# => X"6388d42a",
		16#324c# => X"13860400",
		16#324d# => X"93050000",
		16#324e# => X"13050400",
		16#324f# => X"efa01fa4",
		16#3250# => X"930c0000",
		16#3251# => X"63040500",
		16#3252# => X"b3048540",
		16#3253# => X"138d0c00",
		16#3254# => X"63d49c00",
		16#3255# => X"138d0400",
		16#3256# => X"8346b103",
		16#3257# => X"63840600",
		16#3258# => X"130d1d00",
		16#3259# => X"937d2b00",
		16#325a# => X"63840d00",
		16#325b# => X"130d2d00",
		16#325c# => X"93774b08",
		16#325d# => X"232cf100",
		16#325e# => X"63940706",
		16#325f# => X"b386aa41",
		16#3260# => X"6350d006",
		16#3261# => X"b7470110",
		16#3262# => X"93080001",
		16#3263# => X"1388875e",
		16#3264# => X"13037000",
		16#3265# => X"03264104",
		16#3266# => X"23a00b01",
		16#3267# => X"83258104",
		16#3268# => X"13061600",
		16#3269# => X"13858b00",
		16#326a# => X"63ced848",
		16#326b# => X"23a2db00",
		16#326c# => X"b386b600",
		16#326d# => X"2324d104",
		16#326e# => X"2322c104",
		16#326f# => X"93067000",
		16#3270# => X"930b0500",
		16#3271# => X"63dec600",
		16#3272# => X"13060104",
		16#3273# => X"93050900",
		16#3274# => X"13050a00",
		16#3275# => X"eff0df86",
		16#3276# => X"6312055a",
		16#3277# => X"930bc104",
		16#3278# => X"8346b103",
		16#3279# => X"63880604",
		16#327a# => X"1306b103",
		16#327b# => X"23a0cb00",
		16#327c# => X"13061000",
		16#327d# => X"83264104",
		16#327e# => X"23a2cb00",
		16#327f# => X"03268104",
		16#3280# => X"93861600",
		16#3281# => X"2322d104",
		16#3282# => X"13061600",
		16#3283# => X"2324c104",
		16#3284# => X"13067000",
		16#3285# => X"938b8b00",
		16#3286# => X"635ed600",
		16#3287# => X"13060104",
		16#3288# => X"93050900",
		16#3289# => X"13050a00",
		16#328a# => X"eff09f81",
		16#328b# => X"63180554",
		16#328c# => X"930bc104",
		16#328d# => X"63880d04",
		16#328e# => X"1306c103",
		16#328f# => X"23a0cb00",
		16#3290# => X"13062000",
		16#3291# => X"83264104",
		16#3292# => X"23a2cb00",
		16#3293# => X"03268104",
		16#3294# => X"93861600",
		16#3295# => X"2322d104",
		16#3296# => X"13062600",
		16#3297# => X"2324c104",
		16#3298# => X"13067000",
		16#3299# => X"938b8b00",
		16#329a# => X"635ed600",
		16#329b# => X"13060104",
		16#329c# => X"93050900",
		16#329d# => X"13050a00",
		16#329e# => X"eff08ffc",
		16#329f# => X"63100550",
		16#32a0# => X"930bc104",
		16#32a1# => X"83278101",
		16#32a2# => X"93060008",
		16#32a3# => X"6392d706",
		16#32a4# => X"b38daa41",
		16#32a5# => X"635eb005",
		16#32a6# => X"13080001",
		16#32a7# => X"93087000",
		16#32a8# => X"83270101",
		16#32a9# => X"83264104",
		16#32aa# => X"03268104",
		16#32ab# => X"23a0fb00",
		16#32ac# => X"93861600",
		16#32ad# => X"93858b00",
		16#32ae# => X"6342b83f",
		16#32af# => X"23a2bb01",
		16#32b0# => X"b38dcd00",
		16#32b1# => X"2324b105",
		16#32b2# => X"2322d104",
		16#32b3# => X"13067000",
		16#32b4# => X"938b0500",
		16#32b5# => X"635ed600",
		16#32b6# => X"13060104",
		16#32b7# => X"93050900",
		16#32b8# => X"13050a00",
		16#32b9# => X"eff0cff5",
		16#32ba# => X"631a0548",
		16#32bb# => X"930bc104",
		16#32bc# => X"b38c9c40",
		16#32bd# => X"635e9005",
		16#32be# => X"930d0001",
		16#32bf# => X"13087000",
		16#32c0# => X"83270101",
		16#32c1# => X"83264104",
		16#32c2# => X"03268104",
		16#32c3# => X"23a0fb00",
		16#32c4# => X"93861600",
		16#32c5# => X"93858b00",
		16#32c6# => X"63c69d3d",
		16#32c7# => X"23a29b01",
		16#32c8# => X"b38ccc00",
		16#32c9# => X"23249105",
		16#32ca# => X"2322d104",
		16#32cb# => X"13067000",
		16#32cc# => X"938b0500",
		16#32cd# => X"635ed600",
		16#32ce# => X"13060104",
		16#32cf# => X"93050900",
		16#32d0# => X"13050a00",
		16#32d1# => X"eff0cfef",
		16#32d2# => X"631a0542",
		16#32d3# => X"930bc104",
		16#32d4# => X"83268104",
		16#32d5# => X"23a29b00",
		16#32d6# => X"23a08b00",
		16#32d7# => X"b3849600",
		16#32d8# => X"83264104",
		16#32d9# => X"23249104",
		16#32da# => X"13067000",
		16#32db# => X"93861600",
		16#32dc# => X"2322d104",
		16#32dd# => X"13878b00",
		16#32de# => X"635ed600",
		16#32df# => X"13060104",
		16#32e0# => X"93050900",
		16#32e1# => X"13050a00",
		16#32e2# => X"eff08feb",
		16#32e3# => X"6318053e",
		16#32e4# => X"1307c104",
		16#32e5# => X"93774b00",
		16#32e6# => X"63960738",
		16#32e7# => X"63d4aa01",
		16#32e8# => X"930a0d00",
		16#32e9# => X"83270100",
		16#32ea# => X"b3875701",
		16#32eb# => X"2320f100",
		16#32ec# => X"83278104",
		16#32ed# => X"638c0700",
		16#32ee# => X"13060104",
		16#32ef# => X"93050900",
		16#32f0# => X"13050a00",
		16#32f1# => X"eff0cfe7",
		16#32f2# => X"631a053a",
		16#32f3# => X"23220104",
		16#32f4# => X"130d0c00",
		16#32f5# => X"930bc104",
		16#32f6# => X"6ff0df8f",
		16#32f7# => X"13050400",
		16#32f8# => X"ef405fc3",
		16#32f9# => X"93040500",
		16#32fa# => X"930c0000",
		16#32fb# => X"6ff01fd6",
		16#32fc# => X"136b0b01",
		16#32fd# => X"93760b02",
		16#32fe# => X"63800602",
		16#32ff# => X"130d7d00",
		16#3300# => X"137d8dff",
		16#3301# => X"83280d00",
		16#3302# => X"832c4d00",
		16#3303# => X"130c8d00",
		16#3304# => X"93061000",
		16#3305# => X"6ff05fc7",
		16#3306# => X"93760b01",
		16#3307# => X"130c4d00",
		16#3308# => X"63860600",
		16#3309# => X"83280d00",
		16#330a# => X"6f000001",
		16#330b# => X"93760b04",
		16#330c# => X"63880600",
		16#330d# => X"83580d00",
		16#330e# => X"930c0000",
		16#330f# => X"6ff05ffd",
		16#3310# => X"93760b20",
		16#3311# => X"e38006fe",
		16#3312# => X"83480d00",
		16#3313# => X"6ff0dffe",
		16#3314# => X"b7460110",
		16#3315# => X"93874690",
		16#3316# => X"6ff01f94",
		16#3317# => X"93760b01",
		16#3318# => X"130c4d00",
		16#3319# => X"63860600",
		16#331a# => X"83280d00",
		16#331b# => X"6f000001",
		16#331c# => X"93760b04",
		16#331d# => X"63880600",
		16#331e# => X"83580d00",
		16#331f# => X"930c0000",
		16#3320# => X"6ff09f93",
		16#3321# => X"93760b20",
		16#3322# => X"e38006fe",
		16#3323# => X"83480d00",
		16#3324# => X"6ff0dffe",
		16#3325# => X"13060b00",
		16#3326# => X"93061000",
		16#3327# => X"6ff0dfbf",
		16#3328# => X"13061000",
		16#3329# => X"e38ec6ae",
		16#332a# => X"13062000",
		16#332b# => X"6388c612",
		16#332c# => X"9306010f",
		16#332d# => X"9395dc01",
		16#332e# => X"13f67800",
		16#332f# => X"93d83800",
		16#3330# => X"13060603",
		16#3331# => X"b3e81501",
		16#3332# => X"93dc3c00",
		16#3333# => X"a38fc6fe",
		16#3334# => X"b3e59801",
		16#3335# => X"1384f6ff",
		16#3336# => X"63960502",
		16#3337# => X"93751b00",
		16#3338# => X"638a0500",
		16#3339# => X"93050003",
		16#333a# => X"6306b600",
		16#333b# => X"a30fb4fe",
		16#333c# => X"1384e6ff",
		16#333d# => X"9307010f",
		16#333e# => X"938c0400",
		16#333f# => X"b3848740",
		16#3340# => X"6ff0dfc4",
		16#3341# => X"93060400",
		16#3342# => X"6ff0dffa",
		16#3343# => X"93770b40",
		16#3344# => X"130d0000",
		16#3345# => X"130e010f",
		16#3346# => X"232cf100",
		16#3347# => X"930d9000",
		16#3348# => X"13850800",
		16#3349# => X"1306a000",
		16#334a# => X"93060000",
		16#334b# => X"93850c00",
		16#334c# => X"1304feff",
		16#334d# => X"2322c103",
		16#334e# => X"23201103",
		16#334f# => X"ef005078",
		16#3350# => X"032e4102",
		16#3351# => X"83278101",
		16#3352# => X"13050503",
		16#3353# => X"a30faefe",
		16#3354# => X"130d1d00",
		16#3355# => X"83280102",
		16#3356# => X"638c0704",
		16#3357# => X"83274100",
		16#3358# => X"83c60700",
		16#3359# => X"6396a605",
		16#335a# => X"9307f00f",
		16#335b# => X"6302fd04",
		16#335c# => X"63940c00",
		16#335d# => X"63fe1d03",
		16#335e# => X"8327c100",
		16#335f# => X"83254101",
		16#3360# => X"23201103",
		16#3361# => X"3304f440",
		16#3362# => X"13860700",
		16#3363# => X"13050400",
		16#3364# => X"efc00f82",
		16#3365# => X"83274100",
		16#3366# => X"130d0000",
		16#3367# => X"83280102",
		16#3368# => X"83c61700",
		16#3369# => X"63860600",
		16#336a# => X"93871700",
		16#336b# => X"2322f100",
		16#336c# => X"13850800",
		16#336d# => X"93850c00",
		16#336e# => X"1306a000",
		16#336f# => X"93060000",
		16#3370# => X"ef005012",
		16#3371# => X"938c0500",
		16#3372# => X"b3e5a500",
		16#3373# => X"93080500",
		16#3374# => X"e38205f2",
		16#3375# => X"130e0400",
		16#3376# => X"6ff09ff4",
		16#3377# => X"1304010f",
		16#3378# => X"83278100",
		16#3379# => X"93f6f800",
		16#337a# => X"1304f4ff",
		16#337b# => X"b386d700",
		16#337c# => X"83c60600",
		16#337d# => X"93d84800",
		16#337e# => X"2300d400",
		16#337f# => X"9396cc01",
		16#3380# => X"b3e81601",
		16#3381# => X"93dc4c00",
		16#3382# => X"b3e69801",
		16#3383# => X"e39a06fc",
		16#3384# => X"6ff05fee",
		16#3385# => X"1304010f",
		16#3386# => X"e39e06ec",
		16#3387# => X"13761600",
		16#3388# => X"e30a06ec",
		16#3389# => X"93060003",
		16#338a# => X"a307d10e",
		16#338b# => X"6ff09f98",
		16#338c# => X"63880d1c",
		16#338d# => X"2306b109",
		16#338e# => X"a30d0102",
		16#338f# => X"130c0d00",
		16#3390# => X"6ff0df90",
		16#3391# => X"93850501",
		16#3392# => X"23a21b01",
		16#3393# => X"2324b104",
		16#3394# => X"2322c104",
		16#3395# => X"635ec302",
		16#3396# => X"13060104",
		16#3397# => X"93050900",
		16#3398# => X"13050a00",
		16#3399# => X"23266102",
		16#339a# => X"23240103",
		16#339b# => X"23221103",
		16#339c# => X"2320d102",
		16#339d# => X"eff0cfbc",
		16#339e# => X"63120510",
		16#339f# => X"0323c102",
		16#33a0# => X"03288102",
		16#33a1# => X"83284102",
		16#33a2# => X"83260102",
		16#33a3# => X"1305c104",
		16#33a4# => X"938606ff",
		16#33a5# => X"930b0500",
		16#33a6# => X"6ff0dfaf",
		16#33a7# => X"13060601",
		16#33a8# => X"23a20b01",
		16#33a9# => X"2324c104",
		16#33aa# => X"2322d104",
		16#33ab# => X"63d6d802",
		16#33ac# => X"13060104",
		16#33ad# => X"93050900",
		16#33ae# => X"13050a00",
		16#33af# => X"23201103",
		16#33b0# => X"232c0101",
		16#33b1# => X"eff0cfb7",
		16#33b2# => X"631a050a",
		16#33b3# => X"83280102",
		16#33b4# => X"03288101",
		16#33b5# => X"9305c104",
		16#33b6# => X"938d0dff",
		16#33b7# => X"938b0500",
		16#33b8# => X"6ff01fbc",
		16#33b9# => X"13060601",
		16#33ba# => X"23a2bb01",
		16#33bb# => X"2324c104",
		16#33bc# => X"2322d104",
		16#33bd# => X"6352d802",
		16#33be# => X"13060104",
		16#33bf# => X"93050900",
		16#33c0# => X"13050a00",
		16#33c1# => X"232c0101",
		16#33c2# => X"eff08fb3",
		16#33c3# => X"63180506",
		16#33c4# => X"03288101",
		16#33c5# => X"9305c104",
		16#33c6# => X"938c0cff",
		16#33c7# => X"938b0500",
		16#33c8# => X"6ff01fbe",
		16#33c9# => X"3384aa41",
		16#33ca# => X"e35a80c6",
		16#33cb# => X"b7470110",
		16#33cc# => X"930c0001",
		16#33cd# => X"9384875e",
		16#33ce# => X"930d7000",
		16#33cf# => X"83274104",
		16#33d0# => X"23209700",
		16#33d1# => X"83268104",
		16#33d2# => X"93871700",
		16#33d3# => X"63ce8c06",
		16#33d4# => X"23228700",
		16#33d5# => X"3304d400",
		16#33d6# => X"23248104",
		16#33d7# => X"2322f104",
		16#33d8# => X"13077000",
		16#33d9# => X"e35cf7c2",
		16#33da# => X"13060104",
		16#33db# => X"93050900",
		16#33dc# => X"13050a00",
		16#33dd# => X"eff0cfac",
		16#33de# => X"e30205c2",
		16#33df# => X"8357c900",
		16#33e0# => X"93f70704",
		16#33e1# => X"639e07ce",
		16#33e2# => X"8320c112",
		16#33e3# => X"03248112",
		16#33e4# => X"03250100",
		16#33e5# => X"83244112",
		16#33e6# => X"03290112",
		16#33e7# => X"8329c111",
		16#33e8# => X"032a8111",
		16#33e9# => X"832a4111",
		16#33ea# => X"032b0111",
		16#33eb# => X"832bc110",
		16#33ec# => X"032c8110",
		16#33ed# => X"832c4110",
		16#33ee# => X"032d0110",
		16#33ef# => X"832dc10f",
		16#33f0# => X"13010113",
		16#33f1# => X"67800000",
		16#33f2# => X"93860601",
		16#33f3# => X"23229701",
		16#33f4# => X"2324d104",
		16#33f5# => X"2322f104",
		16#33f6# => X"13078700",
		16#33f7# => X"63defd00",
		16#33f8# => X"13060104",
		16#33f9# => X"93050900",
		16#33fa# => X"13050a00",
		16#33fb# => X"eff04fa5",
		16#33fc# => X"e31605f8",
		16#33fd# => X"1307c104",
		16#33fe# => X"130404ff",
		16#33ff# => X"6ff01ff4",
		16#3400# => X"83278104",
		16#3401# => X"e38c07f6",
		16#3402# => X"13060104",
		16#3403# => X"93050900",
		16#3404# => X"13050a00",
		16#3405# => X"eff0cfa2",
		16#3406# => X"6ff05ff6",
		16#3407# => X"83a7c181",
		16#3408# => X"130101fe",
		16#3409# => X"232c8100",
		16#340a# => X"232a9100",
		16#340b# => X"232e1100",
		16#340c# => X"13040500",
		16#340d# => X"93840600",
		16#340e# => X"83a74703",
		16#340f# => X"63980504",
		16#3410# => X"63960700",
		16#3411# => X"b7570110",
		16#3412# => X"938707ca",
		16#3413# => X"83a7070e",
		16#3414# => X"93860400",
		16#3415# => X"13060000",
		16#3416# => X"93054100",
		16#3417# => X"13050400",
		16#3418# => X"e7800700",
		16#3419# => X"9307f0ff",
		16#341a# => X"6318f500",
		16#341b# => X"23a00400",
		16#341c# => X"9307a008",
		16#341d# => X"2320f400",
		16#341e# => X"8320c101",
		16#341f# => X"03248101",
		16#3420# => X"83244101",
		16#3421# => X"13010102",
		16#3422# => X"67800000",
		16#3423# => X"63960700",
		16#3424# => X"b7570110",
		16#3425# => X"938707ca",
		16#3426# => X"83a7070e",
		16#3427# => X"93860400",
		16#3428# => X"6ff0dffb",
		16#3429# => X"93060600",
		16#342a# => X"13860500",
		16#342b# => X"93050500",
		16#342c# => X"03a5c181",
		16#342d# => X"6ff09ff6",
		16#342e# => X"f32740f1",
		16#342f# => X"b7870110",
		16#3430# => X"37870110",
		16#3431# => X"83a747ab",
		16#3432# => X"032707ab",
		16#3433# => X"13850700",
		16#3434# => X"e7000700",
		16#3435# => X"0b000000",
		16#3436# => X"67800000",
		16#3437# => X"63060500",
		16#3438# => X"0b000000",
		16#3439# => X"6ff0dfff",
		16#343a# => X"67800000",
		16#343b# => X"130101fe",
		16#343c# => X"232c8100",
		16#343d# => X"232a9100",
		16#343e# => X"93040200",
		16#343f# => X"13040200",
		16#3440# => X"23263101",
		16#3441# => X"33848440",
		16#3442# => X"93890500",
		16#3443# => X"b7850110",
		16#3444# => X"23282101",
		16#3445# => X"13060400",
		16#3446# => X"13090500",
		16#3447# => X"938585ab",
		16#3448# => X"13050200",
		16#3449# => X"232e1100",
		16#344a# => X"23244101",
		16#344b# => X"130a0200",
		16#344c# => X"efa00fa7",
		16#344d# => X"13060200",
		16#344e# => X"33069640",
		16#344f# => X"93050000",
		16#3450# => X"33058a00",
		16#3451# => X"efa08fb9",
		16#3452# => X"93850900",
		16#3453# => X"13050900",
		16#3454# => X"eff0dff8",
		16#3455# => X"93050000",
		16#3456# => X"13050000",
		16#3457# => X"ef505020",
		16#3458# => X"ef504061",
		16#3459# => X"130101ff",
		16#345a# => X"23261100",
		16#345b# => X"23248100",
		16#345c# => X"23229100",
		16#345d# => X"732400b0",
		16#345e# => X"f32400b8",
		16#345f# => X"b7c50000",
		16#3460# => X"93850535",
		16#3461# => X"ef50c04a",
		16#3462# => X"b3068500",
		16#3463# => X"33b5a600",
		16#3464# => X"33059500",
		16#3465# => X"732700b0",
		16#3466# => X"f32700b8",
		16#3467# => X"e3eca7fe",
		16#3468# => X"6314f500",
		16#3469# => X"e368d7fe",
		16#346a# => X"8320c100",
		16#346b# => X"03248100",
		16#346c# => X"83244100",
		16#346d# => X"13010101",
		16#346e# => X"67800000",
		16#346f# => X"630c0500",
		16#3470# => X"93071000",
		16#3471# => X"3395a700",
		16#3472# => X"f327207c",
		16#3473# => X"b377f500",
		16#3474# => X"e39c07fe",
		16#3475# => X"63860500",
		16#3476# => X"83a70500",
		16#3477# => X"23a00700",
		16#3478# => X"13050000",
		16#3479# => X"67800000",
		16#347a# => X"130101ff",
		16#347b# => X"23261100",
		16#347c# => X"23248100",
		16#347d# => X"23229100",
		16#347e# => X"23202101",
		16#347f# => X"f328007c",
		16#3480# => X"63eca80a",
		16#3481# => X"635aa00a",
		16#3482# => X"f326107c",
		16#3483# => X"7327207c",
		16#3484# => X"93071000",
		16#3485# => X"9388f8ff",
		16#3486# => X"1305f5ff",
		16#3487# => X"13040000",
		16#3488# => X"63fc1703",
		16#3489# => X"130e1000",
		16#348a# => X"13571700",
		16#348b# => X"93d61600",
		16#348c# => X"13781700",
		16#348d# => X"13f31600",
		16#348e# => X"631c0800",
		16#348f# => X"3318fe00",
		16#3490# => X"63080300",
		16#3491# => X"1305f5ff",
		16#3492# => X"33040401",
		16#3493# => X"63080508",
		16#3494# => X"93871700",
		16#3495# => X"e39af8fc",
		16#3496# => X"63020508",
		16#3497# => X"37450110",
		16#3498# => X"13090600",
		16#3499# => X"93840500",
		16#349a# => X"13860500",
		16#349b# => X"1305059e",
		16#349c# => X"93050400",
		16#349d# => X"ef40cfa4",
		16#349e# => X"b7870110",
		16#349f# => X"23a897aa",
		16#34a0# => X"b7870110",
		16#34a1# => X"23aa27ab",
		16#34a2# => X"b7d70010",
		16#34a3# => X"9387870b",
		16#34a4# => X"93020400",
		16#34a5# => X"13830700",
		16#34a6# => X"8b420300",
		16#34a7# => X"7324247c",
		16#34a8# => X"8320c100",
		16#34a9# => X"03248100",
		16#34aa# => X"83244100",
		16#34ab# => X"03290100",
		16#34ac# => X"13010101",
		16#34ad# => X"67800000",
		16#34ae# => X"03248100",
		16#34af# => X"8320c100",
		16#34b0# => X"83244100",
		16#34b1# => X"03290100",
		16#34b2# => X"93050500",
		16#34b3# => X"37450110",
		16#34b4# => X"13050598",
		16#34b5# => X"13010101",
		16#34b6# => X"6f408f9e",
		16#34b7# => X"03248100",
		16#34b8# => X"8320c100",
		16#34b9# => X"83244100",
		16#34ba# => X"03290100",
		16#34bb# => X"37450110",
		16#34bc# => X"130505a1",
		16#34bd# => X"13010101",
		16#34be# => X"6f404fb9",
		16#34bf# => X"13071000",
		16#34c0# => X"f327207c",
		16#34c1# => X"e39ee7fe",
		16#34c2# => X"67800000",
		16#34c3# => X"130101fe",
		16#34c4# => X"23263101",
		16#34c5# => X"23244101",
		16#34c6# => X"23225101",
		16#34c7# => X"232e1100",
		16#34c8# => X"232c8100",
		16#34c9# => X"232a9100",
		16#34ca# => X"23282101",
		16#34cb# => X"930a0500",
		16#34cc# => X"93890500",
		16#34cd# => X"130a0600",
		16#34ce# => X"7329007c",
		16#34cf# => X"f324107c",
		16#34d0# => X"7324207c",
		16#34d1# => X"37450110",
		16#34d2# => X"13060400",
		16#34d3# => X"93850400",
		16#34d4# => X"130585a4",
		16#34d5# => X"ef40cf96",
		16#34d6# => X"93071000",
		16#34d7# => X"23a00a00",
		16#34d8# => X"63f22703",
		16#34d9# => X"13541400",
		16#34da# => X"93d41400",
		16#34db# => X"13771400",
		16#34dc# => X"93f61400",
		16#34dd# => X"63140700",
		16#34de# => X"63940604",
		16#34df# => X"93871700",
		16#34e0# => X"e312f9fe",
		16#34e1# => X"37450110",
		16#34e2# => X"93850900",
		16#34e3# => X"130505b0",
		16#34e4# => X"ef400f93",
		16#34e5# => X"03248101",
		16#34e6# => X"8320c101",
		16#34e7# => X"83244101",
		16#34e8# => X"03290101",
		16#34e9# => X"832a4100",
		16#34ea# => X"13050a00",
		16#34eb# => X"13830900",
		16#34ec# => X"032a8100",
		16#34ed# => X"8329c100",
		16#34ee# => X"13010102",
		16#34ef# => X"67000300",
		16#34f0# => X"37450110",
		16#34f1# => X"93850700",
		16#34f2# => X"23a0fa00",
		16#34f3# => X"93060a00",
		16#34f4# => X"13860900",
		16#34f5# => X"130585a7",
		16#34f6# => X"13041000",
		16#34f7# => X"3314f400",
		16#34f8# => X"b7840110",
		16#34f9# => X"ef40cf8d",
		16#34fa# => X"37890110",
		16#34fb# => X"03a644ab",
		16#34fc# => X"832509ab",
		16#34fd# => X"b74a0110",
		16#34fe# => X"13854aac",
		16#34ff# => X"ef404f8c",
		16#3500# => X"13060a00",
		16#3501# => X"93850900",
		16#3502# => X"13854aac",
		16#3503# => X"232839ab",
		16#3504# => X"23aa44ab",
		16#3505# => X"ef40cf8a",
		16#3506# => X"b7d70010",
		16#3507# => X"9387870b",
		16#3508# => X"93020400",
		16#3509# => X"13830700",
		16#350a# => X"8b420300",
		16#350b# => X"f327247c",
		16#350c# => X"8320c101",
		16#350d# => X"03248101",
		16#350e# => X"83244101",
		16#350f# => X"03290101",
		16#3510# => X"8329c100",
		16#3511# => X"032a8100",
		16#3512# => X"832a4100",
		16#3513# => X"13010102",
		16#3514# => X"67800000",
		16#3515# => X"67800000",
		16#3516# => X"13051000",
		16#3517# => X"67800000",
		16#3518# => X"130101ff",
		16#3519# => X"23261100",
		16#351a# => X"ef504030",
		16#351b# => X"8320c100",
		16#351c# => X"93076001",
		16#351d# => X"2320f500",
		16#351e# => X"1305f0ff",
		16#351f# => X"13010101",
		16#3520# => X"67800000",
		16#3521# => X"130101ff",
		16#3522# => X"9305f0ff",
		16#3523# => X"23261100",
		16#3524# => X"ef50405b",
		16#3525# => X"0b000000",
		16#3526# => X"6f000000",
		16#3527# => X"6352c004",
		16#3528# => X"03a70183",
		16#3529# => X"9307a000",
		16#352a# => X"03470700",
		16#352b# => X"630af702",
		16#352c# => X"3386c500",
		16#352d# => X"93870500",
		16#352e# => X"1308a000",
		16#352f# => X"6f000001",
		16#3530# => X"03a70183",
		16#3531# => X"03470700",
		16#3532# => X"630e0701",
		16#3533# => X"93871700",
		16#3534# => X"a38fe7fe",
		16#3535# => X"3385b740",
		16#3536# => X"e394c7fe",
		16#3537# => X"67800000",
		16#3538# => X"13050000",
		16#3539# => X"67800000",
		16#353a# => X"83a70183",
		16#353b# => X"2380a700",
		16#353c# => X"67800000",
		16#353d# => X"6352c002",
		16#353e# => X"3388c500",
		16#353f# => X"93851500",
		16#3540# => X"03c7f5ff",
		16#3541# => X"83a70183",
		16#3542# => X"2380e700",
		16#3543# => X"e318b8fe",
		16#3544# => X"13050600",
		16#3545# => X"67800000",
		16#3546# => X"13060000",
		16#3547# => X"13050600",
		16#3548# => X"67800000",
		16#3549# => X"83a78184",
		16#354a# => X"130101ff",
		16#354b# => X"23261100",
		16#354c# => X"63800702",
		16#354d# => X"3385a700",
		16#354e# => X"6364a102",
		16#354f# => X"8320c100",
		16#3550# => X"23a4a184",
		16#3551# => X"13850700",
		16#3552# => X"13010101",
		16#3553# => X"67800000",
		16#3554# => X"93060200",
		16#3555# => X"23a4d184",
		16#3556# => X"93070200",
		16#3557# => X"6ff09ffd",
		16#3558# => X"37450110",
		16#3559# => X"130585b3",
		16#355a# => X"ef404f92",
		16#355b# => X"ef50801e",
		16#355c# => X"1305f0ff",
		16#355d# => X"67800000",
		16#355e# => X"b7270000",
		16#355f# => X"23a2f500",
		16#3560# => X"13050000",
		16#3561# => X"67800000",
		16#3562# => X"13050000",
		16#3563# => X"67800000",
		16#3564# => X"13050000",
		16#3565# => X"67800000",
		16#3566# => X"130101fe",
		16#3567# => X"2324c100",
		16#3568# => X"2326d100",
		16#3569# => X"2328e100",
		16#356a# => X"232af100",
		16#356b# => X"232c0101",
		16#356c# => X"232e1101",
		16#356d# => X"1305f0ff",
		16#356e# => X"13010102",
		16#356f# => X"67800000",
		16#3570# => X"130101ff",
		16#3571# => X"23261100",
		16#3572# => X"ef50401a",
		16#3573# => X"8320c100",
		16#3574# => X"9307a000",
		16#3575# => X"2320f500",
		16#3576# => X"1305f0ff",
		16#3577# => X"13010101",
		16#3578# => X"67800000",
		16#3579# => X"130101ff",
		16#357a# => X"23261100",
		16#357b# => X"ef500018",
		16#357c# => X"8320c100",
		16#357d# => X"93072000",
		16#357e# => X"2320f500",
		16#357f# => X"1305f0ff",
		16#3580# => X"13010101",
		16#3581# => X"67800000",
		16#3582# => X"130101ff",
		16#3583# => X"23248100",
		16#3584# => X"23261100",
		16#3585# => X"23229100",
		16#3586# => X"13040500",
		16#3587# => X"f32400b0",
		16#3588# => X"f32500b8",
		16#3589# => X"37f6fa02",
		16#358a# => X"13850400",
		16#358b# => X"13060608",
		16#358c# => X"93060000",
		16#358d# => X"ef00000b",
		16#358e# => X"2322a400",
		16#358f# => X"2320a400",
		16#3590# => X"2326a400",
		16#3591# => X"2324a400",
		16#3592# => X"8320c100",
		16#3593# => X"03248100",
		16#3594# => X"13850400",
		16#3595# => X"83244100",
		16#3596# => X"13010101",
		16#3597# => X"67800000",
		16#3598# => X"b7270000",
		16#3599# => X"23a2f500",
		16#359a# => X"13050000",
		16#359b# => X"67800000",
		16#359c# => X"130101ff",
		16#359d# => X"23261100",
		16#359e# => X"ef50400f",
		16#359f# => X"8320c100",
		16#35a0# => X"9307f001",
		16#35a1# => X"2320f500",
		16#35a2# => X"1305f0ff",
		16#35a3# => X"13010101",
		16#35a4# => X"67800000",
		16#35a5# => X"130101ff",
		16#35a6# => X"23261100",
		16#35a7# => X"ef50000d",
		16#35a8# => X"8320c100",
		16#35a9# => X"9307b000",
		16#35aa# => X"2320f500",
		16#35ab# => X"1305f0ff",
		16#35ac# => X"13010101",
		16#35ad# => X"67800000",
		16#35ae# => X"130101ff",
		16#35af# => X"23261100",
		16#35b0# => X"ef50c00a",
		16#35b1# => X"8320c100",
		16#35b2# => X"9307c000",
		16#35b3# => X"2320f500",
		16#35b4# => X"1305f0ff",
		16#35b5# => X"13010101",
		16#35b6# => X"67800000",
		16#35b7# => X"13050000",
		16#35b8# => X"67800000",
		16#35b9# => X"130101fd",
		16#35ba# => X"23286101",
		16#35bb# => X"23267101",
		16#35bc# => X"23261102",
		16#35bd# => X"23248102",
		16#35be# => X"23229102",
		16#35bf# => X"23202103",
		16#35c0# => X"232e3101",
		16#35c1# => X"232c4101",
		16#35c2# => X"232a5101",
		16#35c3# => X"23248101",
		16#35c4# => X"23229101",
		16#35c5# => X"2320a101",
		16#35c6# => X"130b0500",
		16#35c7# => X"938b0500",
		16#35c8# => X"639e0638",
		16#35c9# => X"37490110",
		16#35ca# => X"93040600",
		16#35cb# => X"130a0500",
		16#35cc# => X"1309c96b",
		16#35cd# => X"63f8c512",
		16#35ce# => X"b7070100",
		16#35cf# => X"13840500",
		16#35d0# => X"6378f610",
		16#35d1# => X"1307f00f",
		16#35d2# => X"3337c700",
		16#35d3# => X"13173700",
		16#35d4# => X"b357e600",
		16#35d5# => X"3309f900",
		16#35d6# => X"83460900",
		16#35d7# => X"3387e600",
		16#35d8# => X"93060002",
		16#35d9# => X"b386e640",
		16#35da# => X"638c0600",
		16#35db# => X"3394db00",
		16#35dc# => X"3357eb00",
		16#35dd# => X"b314d600",
		16#35de# => X"33648700",
		16#35df# => X"331adb00",
		16#35e0# => X"93da0401",
		16#35e1# => X"93850a00",
		16#35e2# => X"13050400",
		16#35e3# => X"ef409071",
		16#35e4# => X"93090500",
		16#35e5# => X"93850a00",
		16#35e6# => X"13050400",
		16#35e7# => X"139b0401",
		16#35e8# => X"ef40d06b",
		16#35e9# => X"135b0b01",
		16#35ea# => X"13090500",
		16#35eb# => X"93050500",
		16#35ec# => X"13050b00",
		16#35ed# => X"ef40d067",
		16#35ee# => X"93990901",
		16#35ef# => X"93570a01",
		16#35f0# => X"b3e7f900",
		16#35f1# => X"13040900",
		16#35f2# => X"63fea700",
		16#35f3# => X"b3879700",
		16#35f4# => X"1304f9ff",
		16#35f5# => X"63e89700",
		16#35f6# => X"63f6a700",
		16#35f7# => X"1304e9ff",
		16#35f8# => X"b3879700",
		16#35f9# => X"3389a740",
		16#35fa# => X"93850a00",
		16#35fb# => X"13050900",
		16#35fc# => X"ef40506b",
		16#35fd# => X"93090500",
		16#35fe# => X"93850a00",
		16#35ff# => X"13050900",
		16#3600# => X"ef40d065",
		16#3601# => X"131a0a01",
		16#3602# => X"13090500",
		16#3603# => X"93050500",
		16#3604# => X"93990901",
		16#3605# => X"13050b00",
		16#3606# => X"135a0a01",
		16#3607# => X"ef405061",
		16#3608# => X"33ea4901",
		16#3609# => X"13060900",
		16#360a# => X"637caa00",
		16#360b# => X"338a4401",
		16#360c# => X"1306f9ff",
		16#360d# => X"63669a00",
		16#360e# => X"6374aa00",
		16#360f# => X"1306e9ff",
		16#3610# => X"13140401",
		16#3611# => X"3364c400",
		16#3612# => X"930a0000",
		16#3613# => X"6f000013",
		16#3614# => X"b7070001",
		16#3615# => X"13070001",
		16#3616# => X"e36cf6ee",
		16#3617# => X"13078001",
		16#3618# => X"6ff01fef",
		16#3619# => X"93890600",
		16#361a# => X"631a0600",
		16#361b# => X"93050000",
		16#361c# => X"13051000",
		16#361d# => X"ef40905e",
		16#361e# => X"93040500",
		16#361f# => X"b7070100",
		16#3620# => X"63fef412",
		16#3621# => X"9307f00f",
		16#3622# => X"63f49700",
		16#3623# => X"93098000",
		16#3624# => X"b3d73401",
		16#3625# => X"3309f900",
		16#3626# => X"03470900",
		16#3627# => X"93060002",
		16#3628# => X"33073701",
		16#3629# => X"b386e640",
		16#362a# => X"63940612",
		16#362b# => X"33849b40",
		16#362c# => X"930a1000",
		16#362d# => X"13db0401",
		16#362e# => X"93050b00",
		16#362f# => X"13050400",
		16#3630# => X"ef40505e",
		16#3631# => X"93090500",
		16#3632# => X"93050b00",
		16#3633# => X"13050400",
		16#3634# => X"939b0401",
		16#3635# => X"ef409058",
		16#3636# => X"93db0b01",
		16#3637# => X"13090500",
		16#3638# => X"93050500",
		16#3639# => X"13850b00",
		16#363a# => X"ef409054",
		16#363b# => X"93990901",
		16#363c# => X"93570a01",
		16#363d# => X"b3e7f900",
		16#363e# => X"13040900",
		16#363f# => X"63fea700",
		16#3640# => X"b3879700",
		16#3641# => X"1304f9ff",
		16#3642# => X"63e89700",
		16#3643# => X"63f6a700",
		16#3644# => X"1304e9ff",
		16#3645# => X"b3879700",
		16#3646# => X"3389a740",
		16#3647# => X"93050b00",
		16#3648# => X"13050900",
		16#3649# => X"ef401058",
		16#364a# => X"93090500",
		16#364b# => X"93050b00",
		16#364c# => X"13050900",
		16#364d# => X"ef409052",
		16#364e# => X"131a0a01",
		16#364f# => X"13090500",
		16#3650# => X"93050500",
		16#3651# => X"93990901",
		16#3652# => X"13850b00",
		16#3653# => X"135a0a01",
		16#3654# => X"ef40104e",
		16#3655# => X"33ea4901",
		16#3656# => X"13060900",
		16#3657# => X"637caa00",
		16#3658# => X"338a4401",
		16#3659# => X"1306f9ff",
		16#365a# => X"63669a00",
		16#365b# => X"6374aa00",
		16#365c# => X"1306e9ff",
		16#365d# => X"13140401",
		16#365e# => X"3364c400",
		16#365f# => X"13050400",
		16#3660# => X"93850a00",
		16#3661# => X"8320c102",
		16#3662# => X"03248102",
		16#3663# => X"83244102",
		16#3664# => X"03290102",
		16#3665# => X"8329c101",
		16#3666# => X"032a8101",
		16#3667# => X"832a4101",
		16#3668# => X"032b0101",
		16#3669# => X"832bc100",
		16#366a# => X"032c8100",
		16#366b# => X"832c4100",
		16#366c# => X"032d0100",
		16#366d# => X"13010103",
		16#366e# => X"67800000",
		16#366f# => X"b7070001",
		16#3670# => X"93090001",
		16#3671# => X"e3e6f4ec",
		16#3672# => X"93098001",
		16#3673# => X"6ff05fec",
		16#3674# => X"b394d400",
		16#3675# => X"b3d9eb00",
		16#3676# => X"13d40401",
		16#3677# => X"3357eb00",
		16#3678# => X"b39bdb00",
		16#3679# => X"93050400",
		16#367a# => X"13850900",
		16#367b# => X"b36b7701",
		16#367c# => X"331adb00",
		16#367d# => X"ef40104b",
		16#367e# => X"13090500",
		16#367f# => X"93050400",
		16#3680# => X"13850900",
		16#3681# => X"139b0401",
		16#3682# => X"ef405045",
		16#3683# => X"135b0b01",
		16#3684# => X"93090500",
		16#3685# => X"93050500",
		16#3686# => X"13050b00",
		16#3687# => X"ef405041",
		16#3688# => X"13190901",
		16#3689# => X"13d70b01",
		16#368a# => X"3367e900",
		16#368b# => X"938a0900",
		16#368c# => X"637ea700",
		16#368d# => X"33079700",
		16#368e# => X"938af9ff",
		16#368f# => X"63689700",
		16#3690# => X"6376a700",
		16#3691# => X"938ae9ff",
		16#3692# => X"33079700",
		16#3693# => X"b309a740",
		16#3694# => X"93050400",
		16#3695# => X"13850900",
		16#3696# => X"ef40d044",
		16#3697# => X"93050400",
		16#3698# => X"13090500",
		16#3699# => X"13850900",
		16#369a# => X"ef40503f",
		16#369b# => X"13040500",
		16#369c# => X"93050500",
		16#369d# => X"13050b00",
		16#369e# => X"ef40903b",
		16#369f# => X"13970b01",
		16#36a0# => X"13570701",
		16#36a1# => X"13190901",
		16#36a2# => X"b367e900",
		16#36a3# => X"13070400",
		16#36a4# => X"63fea700",
		16#36a5# => X"b3879700",
		16#36a6# => X"1307f4ff",
		16#36a7# => X"63e89700",
		16#36a8# => X"63f6a700",
		16#36a9# => X"1307e4ff",
		16#36aa# => X"b3879700",
		16#36ab# => X"939a0a01",
		16#36ac# => X"3384a740",
		16#36ad# => X"b3eaea00",
		16#36ae# => X"6ff0dfdf",
		16#36af# => X"63ecd51e",
		16#36b0# => X"b7070100",
		16#36b1# => X"63f4f604",
		16#36b2# => X"1307f00f",
		16#36b3# => X"b335d700",
		16#36b4# => X"93953500",
		16#36b5# => X"37470110",
		16#36b6# => X"1307c76b",
		16#36b7# => X"b3d7b600",
		16#36b8# => X"b387e700",
		16#36b9# => X"03c70700",
		16#36ba# => X"930a0002",
		16#36bb# => X"3307b700",
		16#36bc# => X"b38aea40",
		16#36bd# => X"63960a02",
		16#36be# => X"13041000",
		16#36bf# => X"e3e076e9",
		16#36c0# => X"3336cb00",
		16#36c1# => X"13441600",
		16#36c2# => X"6ff05fe7",
		16#36c3# => X"b7070001",
		16#36c4# => X"93050001",
		16#36c5# => X"e3e0f6fc",
		16#36c6# => X"93058001",
		16#36c7# => X"6ff09ffb",
		16#36c8# => X"b35ce600",
		16#36c9# => X"b3965601",
		16#36ca# => X"b3ecdc00",
		16#36cb# => X"b3d4eb00",
		16#36cc# => X"b3975b01",
		16#36cd# => X"93db0c01",
		16#36ce# => X"3357eb00",
		16#36cf# => X"93850b00",
		16#36d0# => X"13850400",
		16#36d1# => X"3364f700",
		16#36d2# => X"b3195601",
		16#36d3# => X"ef409035",
		16#36d4# => X"13090500",
		16#36d5# => X"93850b00",
		16#36d6# => X"13850400",
		16#36d7# => X"139c0c01",
		16#36d8# => X"ef40d02f",
		16#36d9# => X"135c0c01",
		16#36da# => X"93040500",
		16#36db# => X"93050500",
		16#36dc# => X"13050c00",
		16#36dd# => X"ef40d02b",
		16#36de# => X"13190901",
		16#36df# => X"13570401",
		16#36e0# => X"3367e900",
		16#36e1# => X"138a0400",
		16#36e2# => X"637ea700",
		16#36e3# => X"33079701",
		16#36e4# => X"138af4ff",
		16#36e5# => X"63689701",
		16#36e6# => X"6376a700",
		16#36e7# => X"138ae4ff",
		16#36e8# => X"33079701",
		16#36e9# => X"b304a740",
		16#36ea# => X"93850b00",
		16#36eb# => X"13850400",
		16#36ec# => X"ef40502f",
		16#36ed# => X"13090500",
		16#36ee# => X"93850b00",
		16#36ef# => X"13850400",
		16#36f0# => X"ef40d029",
		16#36f1# => X"93040500",
		16#36f2# => X"93050500",
		16#36f3# => X"13050c00",
		16#36f4# => X"ef401026",
		16#36f5# => X"93170401",
		16#36f6# => X"13190901",
		16#36f7# => X"93d70701",
		16#36f8# => X"b367f900",
		16#36f9# => X"13860400",
		16#36fa# => X"63fea700",
		16#36fb# => X"b3879701",
		16#36fc# => X"1386f4ff",
		16#36fd# => X"63e89701",
		16#36fe# => X"63f6a700",
		16#36ff# => X"1386e4ff",
		16#3700# => X"b3879701",
		16#3701# => X"13140a01",
		16#3702# => X"b70b0100",
		16#3703# => X"3364c400",
		16#3704# => X"1389fbff",
		16#3705# => X"337d2401",
		16#3706# => X"33f92901",
		16#3707# => X"b384a740",
		16#3708# => X"93050900",
		16#3709# => X"13050d00",
		16#370a# => X"ef409020",
		16#370b# => X"935c0401",
		16#370c# => X"93050900",
		16#370d# => X"130a0500",
		16#370e# => X"13850c00",
		16#370f# => X"ef40501f",
		16#3710# => X"93d90901",
		16#3711# => X"130c0500",
		16#3712# => X"93850900",
		16#3713# => X"13850c00",
		16#3714# => X"ef40101e",
		16#3715# => X"13090500",
		16#3716# => X"93850900",
		16#3717# => X"13050d00",
		16#3718# => X"ef40101d",
		16#3719# => X"33058501",
		16#371a# => X"93570a01",
		16#371b# => X"3385a700",
		16#371c# => X"63748501",
		16#371d# => X"33097901",
		16#371e# => X"93570501",
		16#371f# => X"b3872701",
		16#3720# => X"63e6f402",
		16#3721# => X"e392f4bc",
		16#3722# => X"b7070100",
		16#3723# => X"9387f7ff",
		16#3724# => X"3375f500",
		16#3725# => X"13150501",
		16#3726# => X"337afa00",
		16#3727# => X"33165b01",
		16#3728# => X"33054501",
		16#3729# => X"930a0000",
		16#372a# => X"e37aa6cc",
		16#372b# => X"1304f4ff",
		16#372c# => X"6ff09fb9",
		16#372d# => X"930a0000",
		16#372e# => X"13040000",
		16#372f# => X"6ff01fcc",
		16#3730# => X"130101fb",
		16#3731# => X"23248104",
		16#3732# => X"23229104",
		16#3733# => X"232e3103",
		16#3734# => X"23229103",
		16#3735# => X"23261104",
		16#3736# => X"23202105",
		16#3737# => X"232c4103",
		16#3738# => X"232a5103",
		16#3739# => X"23286103",
		16#373a# => X"23267103",
		16#373b# => X"23248103",
		16#373c# => X"2320a103",
		16#373d# => X"232eb101",
		16#373e# => X"930c0500",
		16#373f# => X"93890500",
		16#3740# => X"13040500",
		16#3741# => X"93840500",
		16#3742# => X"639e0626",
		16#3743# => X"b74a0110",
		16#3744# => X"13090600",
		16#3745# => X"138a0600",
		16#3746# => X"938aca6b",
		16#3747# => X"63f4c514",
		16#3748# => X"b7070100",
		16#3749# => X"6376f612",
		16#374a# => X"9307f00f",
		16#374b# => X"63f4c700",
		16#374c# => X"130a8000",
		16#374d# => X"b3574601",
		16#374e# => X"b38afa00",
		16#374f# => X"03c70a00",
		16#3750# => X"13050002",
		16#3751# => X"33074701",
		16#3752# => X"330ae540",
		16#3753# => X"630c0a00",
		16#3754# => X"b3954901",
		16#3755# => X"33d7ec00",
		16#3756# => X"33194601",
		16#3757# => X"b364b700",
		16#3758# => X"33944c01",
		16#3759# => X"935a0901",
		16#375a# => X"93850a00",
		16#375b# => X"13850400",
		16#375c# => X"ef405013",
		16#375d# => X"93090500",
		16#375e# => X"93850a00",
		16#375f# => X"131b0901",
		16#3760# => X"13850400",
		16#3761# => X"ef40900d",
		16#3762# => X"135b0b01",
		16#3763# => X"93050500",
		16#3764# => X"13050b00",
		16#3765# => X"ef40d009",
		16#3766# => X"93990901",
		16#3767# => X"93570401",
		16#3768# => X"b3e7f900",
		16#3769# => X"63faa700",
		16#376a# => X"b3872701",
		16#376b# => X"63e62701",
		16#376c# => X"63f4a700",
		16#376d# => X"b3872701",
		16#376e# => X"b384a740",
		16#376f# => X"93850a00",
		16#3770# => X"13850400",
		16#3771# => X"ef40100e",
		16#3772# => X"93090500",
		16#3773# => X"93850a00",
		16#3774# => X"13850400",
		16#3775# => X"ef409008",
		16#3776# => X"13140401",
		16#3777# => X"93050500",
		16#3778# => X"93990901",
		16#3779# => X"13050b00",
		16#377a# => X"13540401",
		16#377b# => X"ef405004",
		16#377c# => X"33e48900",
		16#377d# => X"637aa400",
		16#377e# => X"33042401",
		16#377f# => X"63662401",
		16#3780# => X"6374a400",
		16#3781# => X"33042401",
		16#3782# => X"3304a440",
		16#3783# => X"33554401",
		16#3784# => X"93050000",
		16#3785# => X"8320c104",
		16#3786# => X"03248104",
		16#3787# => X"83244104",
		16#3788# => X"03290104",
		16#3789# => X"8329c103",
		16#378a# => X"032a8103",
		16#378b# => X"832a4103",
		16#378c# => X"032b0103",
		16#378d# => X"832bc102",
		16#378e# => X"032c8102",
		16#378f# => X"832c4102",
		16#3790# => X"032d0102",
		16#3791# => X"832dc101",
		16#3792# => X"13010105",
		16#3793# => X"67800000",
		16#3794# => X"b7070001",
		16#3795# => X"130a0001",
		16#3796# => X"e36ef6ec",
		16#3797# => X"130a8001",
		16#3798# => X"6ff05fed",
		16#3799# => X"631a0600",
		16#379a# => X"93050000",
		16#379b# => X"13051000",
		16#379c# => X"ef40c07e",
		16#379d# => X"13090500",
		16#379e# => X"b7070100",
		16#379f# => X"637af90e",
		16#37a0# => X"9307f00f",
		16#37a1# => X"63f42701",
		16#37a2# => X"130a8000",
		16#37a3# => X"b3574901",
		16#37a4# => X"b38afa00",
		16#37a5# => X"03c70a00",
		16#37a6# => X"13050002",
		16#37a7# => X"b3842941",
		16#37a8# => X"33074701",
		16#37a9# => X"330ae540",
		16#37aa# => X"e30e0aea",
		16#37ab# => X"33194901",
		16#37ac# => X"b3dae900",
		16#37ad# => X"b3954901",
		16#37ae# => X"33d7ec00",
		16#37af# => X"93540901",
		16#37b0# => X"336bb700",
		16#37b1# => X"13850a00",
		16#37b2# => X"93850400",
		16#37b3# => X"ef40807d",
		16#37b4# => X"93090500",
		16#37b5# => X"93850400",
		16#37b6# => X"931b0901",
		16#37b7# => X"13850a00",
		16#37b8# => X"ef40c077",
		16#37b9# => X"93db0b01",
		16#37ba# => X"93050500",
		16#37bb# => X"13850b00",
		16#37bc# => X"ef400074",
		16#37bd# => X"93990901",
		16#37be# => X"93570b01",
		16#37bf# => X"b3e7f900",
		16#37c0# => X"33944c01",
		16#37c1# => X"63faa700",
		16#37c2# => X"b3872701",
		16#37c3# => X"63e62701",
		16#37c4# => X"63f4a700",
		16#37c5# => X"b3872701",
		16#37c6# => X"b38aa740",
		16#37c7# => X"93850400",
		16#37c8# => X"13850a00",
		16#37c9# => X"ef400078",
		16#37ca# => X"93090500",
		16#37cb# => X"93850400",
		16#37cc# => X"13850a00",
		16#37cd# => X"ef408072",
		16#37ce# => X"93050500",
		16#37cf# => X"13850b00",
		16#37d0# => X"ef40006f",
		16#37d1# => X"93150b01",
		16#37d2# => X"93990901",
		16#37d3# => X"93d50501",
		16#37d4# => X"b3e5b900",
		16#37d5# => X"63faa500",
		16#37d6# => X"b3852501",
		16#37d7# => X"63e62501",
		16#37d8# => X"63f4a500",
		16#37d9# => X"b3852501",
		16#37da# => X"b384a540",
		16#37db# => X"6ff09fdf",
		16#37dc# => X"b7070001",
		16#37dd# => X"130a0001",
		16#37de# => X"e36af9f0",
		16#37df# => X"130a8001",
		16#37e0# => X"6ff0dff0",
		16#37e1# => X"e3e8d5e8",
		16#37e2# => X"b7070100",
		16#37e3# => X"63fcf604",
		16#37e4# => X"930bf00f",
		16#37e5# => X"33b5db00",
		16#37e6# => X"13153500",
		16#37e7# => X"37470110",
		16#37e8# => X"b3d7a600",
		16#37e9# => X"1307c76b",
		16#37ea# => X"b387e700",
		16#37eb# => X"83cb0700",
		16#37ec# => X"93050002",
		16#37ed# => X"b38bab00",
		16#37ee# => X"338b7541",
		16#37ef# => X"631e0b02",
		16#37f0# => X"63e43601",
		16#37f1# => X"63eacc00",
		16#37f2# => X"3384cc40",
		16#37f3# => X"b386d940",
		16#37f4# => X"33b58c00",
		16#37f5# => X"b384a640",
		16#37f6# => X"13050400",
		16#37f7# => X"93850400",
		16#37f8# => X"6ff05fe3",
		16#37f9# => X"b7070001",
		16#37fa# => X"13050001",
		16#37fb# => X"e3e8f6fa",
		16#37fc# => X"13058001",
		16#37fd# => X"6ff09ffa",
		16#37fe# => X"b3966601",
		16#37ff# => X"335d7601",
		16#3800# => X"336ddd00",
		16#3801# => X"33d47901",
		16#3802# => X"b3956901",
		16#3803# => X"33dc7c01",
		16#3804# => X"93540d01",
		16#3805# => X"336cbc00",
		16#3806# => X"13050400",
		16#3807# => X"93850400",
		16#3808# => X"b31a6601",
		16#3809# => X"ef400068",
		16#380a# => X"130a0500",
		16#380b# => X"93850400",
		16#380c# => X"13050400",
		16#380d# => X"33996c01",
		16#380e# => X"931c0d01",
		16#380f# => X"ef400062",
		16#3810# => X"93dc0c01",
		16#3811# => X"13040500",
		16#3812# => X"93050500",
		16#3813# => X"13850c00",
		16#3814# => X"ef40005e",
		16#3815# => X"131a0a01",
		16#3816# => X"13570c01",
		16#3817# => X"3367ea00",
		16#3818# => X"130a0400",
		16#3819# => X"637ea700",
		16#381a# => X"3307a701",
		16#381b# => X"130af4ff",
		16#381c# => X"6368a701",
		16#381d# => X"6376a700",
		16#381e# => X"130ae4ff",
		16#381f# => X"3307a701",
		16#3820# => X"b309a740",
		16#3821# => X"93850400",
		16#3822# => X"13850900",
		16#3823# => X"ef408061",
		16#3824# => X"93850400",
		16#3825# => X"13040500",
		16#3826# => X"13850900",
		16#3827# => X"ef40005c",
		16#3828# => X"93050500",
		16#3829# => X"93040500",
		16#382a# => X"13850c00",
		16#382b# => X"ef404058",
		16#382c# => X"93150c01",
		16#382d# => X"13140401",
		16#382e# => X"93d50501",
		16#382f# => X"b365b400",
		16#3830# => X"13870400",
		16#3831# => X"63fea500",
		16#3832# => X"b385a501",
		16#3833# => X"1387f4ff",
		16#3834# => X"63e8a501",
		16#3835# => X"63f6a500",
		16#3836# => X"1387e4ff",
		16#3837# => X"b385a501",
		16#3838# => X"131a0a01",
		16#3839# => X"b70c0100",
		16#383a# => X"336aea00",
		16#383b# => X"1384fcff",
		16#383c# => X"b3778a00",
		16#383d# => X"33f48a00",
		16#383e# => X"b384a540",
		16#383f# => X"13850700",
		16#3840# => X"93050400",
		16#3841# => X"2326f100",
		16#3842# => X"135a0a01",
		16#3843# => X"ef404052",
		16#3844# => X"93090500",
		16#3845# => X"93050400",
		16#3846# => X"13050a00",
		16#3847# => X"ef404051",
		16#3848# => X"13dc0a01",
		16#3849# => X"930d0500",
		16#384a# => X"93050c00",
		16#384b# => X"13050a00",
		16#384c# => X"ef400050",
		16#384d# => X"8327c100",
		16#384e# => X"130a0500",
		16#384f# => X"93050c00",
		16#3850# => X"13850700",
		16#3851# => X"ef40c04e",
		16#3852# => X"3305b501",
		16#3853# => X"13d70901",
		16#3854# => X"3307a700",
		16#3855# => X"6374b701",
		16#3856# => X"330a9a01",
		16#3857# => X"b7070100",
		16#3858# => X"9387f7ff",
		16#3859# => X"93550701",
		16#385a# => X"3377f700",
		16#385b# => X"13170701",
		16#385c# => X"b3f7f900",
		16#385d# => X"b3854501",
		16#385e# => X"b307f700",
		16#385f# => X"63e6b400",
		16#3860# => X"639eb400",
		16#3861# => X"637cf900",
		16#3862# => X"33865741",
		16#3863# => X"b3b7c700",
		16#3864# => X"b385a541",
		16#3865# => X"b385f540",
		16#3866# => X"93070600",
		16#3867# => X"b307f940",
		16#3868# => X"3339f900",
		16#3869# => X"b385b440",
		16#386a# => X"b3852541",
		16#386b# => X"33947501",
		16#386c# => X"b3d76701",
		16#386d# => X"3365f400",
		16#386e# => X"b3d56501",
		16#386f# => X"6ff09fc5",
		16#3870# => X"130101fb",
		16#3871# => X"23248104",
		16#3872# => X"232c4103",
		16#3873# => X"37041000",
		16#3874# => X"13da4501",
		16#3875# => X"23202105",
		16#3876# => X"232e3103",
		16#3877# => X"232a5103",
		16#3878# => X"23248103",
		16#3879# => X"1304f4ff",
		16#387a# => X"23261104",
		16#387b# => X"23229104",
		16#387c# => X"23286103",
		16#387d# => X"23267103",
		16#387e# => X"23229103",
		16#387f# => X"2320a103",
		16#3880# => X"232eb101",
		16#3881# => X"137afa7f",
		16#3882# => X"13090500",
		16#3883# => X"130c0600",
		16#3884# => X"938a0600",
		16#3885# => X"3374b400",
		16#3886# => X"93d9f501",
		16#3887# => X"63040a0a",
		16#3888# => X"9307f07f",
		16#3889# => X"6302fa10",
		16#388a# => X"13143400",
		16#388b# => X"b7078000",
		16#388c# => X"3364f400",
		16#388d# => X"135bd501",
		16#388e# => X"336b8b00",
		16#388f# => X"93143500",
		16#3890# => X"130a1ac0",
		16#3891# => X"930b0000",
		16#3892# => X"13d54a01",
		16#3893# => X"37091000",
		16#3894# => X"1309f9ff",
		16#3895# => X"1375f57f",
		16#3896# => X"33795901",
		16#3897# => X"93050c00",
		16#3898# => X"93dafa01",
		16#3899# => X"63000510",
		16#389a# => X"9307f07f",
		16#389b# => X"6300f516",
		16#389c# => X"37048000",
		16#389d# => X"13193900",
		16#389e# => X"33698900",
		16#389f# => X"1354dc01",
		16#38a0# => X"33642401",
		16#38a1# => X"93153c00",
		16#38a2# => X"130515c0",
		16#38a3# => X"93070000",
		16#38a4# => X"13972b00",
		16#38a5# => X"3367f700",
		16#38a6# => X"1307f7ff",
		16#38a7# => X"9306e000",
		16#38a8# => X"33c95901",
		16#38a9# => X"330aaa40",
		16#38aa# => X"63eee614",
		16#38ab# => X"b7460110",
		16#38ac# => X"13172700",
		16#38ad# => X"93868660",
		16#38ae# => X"3307d700",
		16#38af# => X"03270700",
		16#38b0# => X"67000700",
		16#38b1# => X"336ba400",
		16#38b2# => X"630e0b06",
		16#38b3# => X"63000404",
		16#38b4# => X"13050400",
		16#38b5# => X"ef404043",
		16#38b6# => X"930755ff",
		16#38b7# => X"1307c001",
		16#38b8# => X"634cf702",
		16#38b9# => X"130bd001",
		16#38ba# => X"930485ff",
		16#38bb# => X"330bfb40",
		16#38bc# => X"33149400",
		16#38bd# => X"335b6901",
		16#38be# => X"336b8b00",
		16#38bf# => X"b3149900",
		16#38c0# => X"130ad0c0",
		16#38c1# => X"330aaa40",
		16#38c2# => X"6ff0dff3",
		16#38c3# => X"ef40c03f",
		16#38c4# => X"13050502",
		16#38c5# => X"6ff05ffc",
		16#38c6# => X"130485fd",
		16#38c7# => X"331b8900",
		16#38c8# => X"93040000",
		16#38c9# => X"6ff0dffd",
		16#38ca# => X"336ba400",
		16#38cb# => X"63040b02",
		16#38cc# => X"93040500",
		16#38cd# => X"130b0400",
		16#38ce# => X"130af07f",
		16#38cf# => X"930b3000",
		16#38d0# => X"6ff09ff0",
		16#38d1# => X"93040000",
		16#38d2# => X"130a0000",
		16#38d3# => X"930b1000",
		16#38d4# => X"6ff09fef",
		16#38d5# => X"93040000",
		16#38d6# => X"130af07f",
		16#38d7# => X"930b2000",
		16#38d8# => X"6ff09fee",
		16#38d9# => X"33648901",
		16#38da# => X"630e0406",
		16#38db# => X"63000904",
		16#38dc# => X"13050900",
		16#38dd# => X"ef404039",
		16#38de# => X"930755ff",
		16#38df# => X"1307c001",
		16#38e0# => X"634ef702",
		16#38e1# => X"1304d001",
		16#38e2# => X"930585ff",
		16#38e3# => X"3304f440",
		16#38e4# => X"3319b900",
		16#38e5# => X"33548c00",
		16#38e6# => X"33642401",
		16#38e7# => X"b315bc00",
		16#38e8# => X"1307d0c0",
		16#38e9# => X"3305a740",
		16#38ea# => X"6ff05fee",
		16#38eb# => X"13050c00",
		16#38ec# => X"ef408035",
		16#38ed# => X"13050502",
		16#38ee# => X"6ff01ffc",
		16#38ef# => X"130485fd",
		16#38f0# => X"33148c00",
		16#38f1# => X"93050000",
		16#38f2# => X"6ff09ffd",
		16#38f3# => X"33648901",
		16#38f4# => X"63020402",
		16#38f5# => X"13040900",
		16#38f6# => X"1305f07f",
		16#38f7# => X"93073000",
		16#38f8# => X"6ff01feb",
		16#38f9# => X"93050000",
		16#38fa# => X"13050000",
		16#38fb# => X"93071000",
		16#38fc# => X"6ff01fea",
		16#38fd# => X"93050000",
		16#38fe# => X"1305f07f",
		16#38ff# => X"93072000",
		16#3900# => X"6ff01fe9",
		16#3901# => X"63666401",
		16#3902# => X"63128b48",
		16#3903# => X"63e0b448",
		16#3904# => X"9316fb01",
		16#3905# => X"13d71400",
		16#3906# => X"139cf401",
		16#3907# => X"135b1b00",
		16#3908# => X"b3e4e600",
		16#3909# => X"13148400",
		16#390a# => X"93dc8501",
		16#390b# => X"b3ec8c00",
		16#390c# => X"93da0c01",
		16#390d# => X"93970c01",
		16#390e# => X"93d70701",
		16#390f# => X"139d8500",
		16#3910# => X"13050b00",
		16#3911# => X"93850a00",
		16#3912# => X"2322f100",
		16#3913# => X"ef400021",
		16#3914# => X"93050500",
		16#3915# => X"930b0500",
		16#3916# => X"13950c01",
		16#3917# => X"13550501",
		16#3918# => X"ef40001d",
		16#3919# => X"13040500",
		16#391a# => X"93850a00",
		16#391b# => X"13050b00",
		16#391c# => X"ef404023",
		16#391d# => X"13150501",
		16#391e# => X"13d70401",
		16#391f# => X"3365a700",
		16#3920# => X"93890b00",
		16#3921# => X"637e8500",
		16#3922# => X"33059501",
		16#3923# => X"9389fbff",
		16#3924# => X"63689501",
		16#3925# => X"63768500",
		16#3926# => X"9389ebff",
		16#3927# => X"33059501",
		16#3928# => X"33048540",
		16#3929# => X"93850a00",
		16#392a# => X"13050400",
		16#392b# => X"ef40001b",
		16#392c# => X"93050500",
		16#392d# => X"930b0500",
		16#392e# => X"13950c01",
		16#392f# => X"13550501",
		16#3930# => X"ef400017",
		16#3931# => X"130b0500",
		16#3932# => X"93850a00",
		16#3933# => X"13050400",
		16#3934# => X"ef40401d",
		16#3935# => X"939d0401",
		16#3936# => X"13150501",
		16#3937# => X"93dd0d01",
		16#3938# => X"b3edad00",
		16#3939# => X"13870b00",
		16#393a# => X"63fe6d01",
		16#393b# => X"b38d9d01",
		16#393c# => X"1387fbff",
		16#393d# => X"63e89d01",
		16#393e# => X"63f66d01",
		16#393f# => X"1387ebff",
		16#3940# => X"b38d9d01",
		16#3941# => X"93960901",
		16#3942# => X"b7040100",
		16#3943# => X"b3e6e600",
		16#3944# => X"b38d6d41",
		16#3945# => X"138bf4ff",
		16#3946# => X"33f76601",
		16#3947# => X"337b6d01",
		16#3948# => X"13050700",
		16#3949# => X"93050b00",
		16#394a# => X"13d40601",
		16#394b# => X"2326d100",
		16#394c# => X"2324e100",
		16#394d# => X"ef40c00f",
		16#394e# => X"2322a100",
		16#394f# => X"93050b00",
		16#3950# => X"13050400",
		16#3951# => X"ef40c00e",
		16#3952# => X"935b0d01",
		16#3953# => X"93090500",
		16#3954# => X"93850b00",
		16#3955# => X"13050400",
		16#3956# => X"ef40800d",
		16#3957# => X"03278100",
		16#3958# => X"13040500",
		16#3959# => X"13850b00",
		16#395a# => X"93050700",
		16#395b# => X"ef40400c",
		16#395c# => X"03264100",
		16#395d# => X"33053501",
		16#395e# => X"8326c100",
		16#395f# => X"13570601",
		16#3960# => X"3307a700",
		16#3961# => X"63743701",
		16#3962# => X"33049400",
		16#3963# => X"37050100",
		16#3964# => X"1305f5ff",
		16#3965# => X"93540701",
		16#3966# => X"b379a700",
		16#3967# => X"93990901",
		16#3968# => X"3376a600",
		16#3969# => X"b3848400",
		16#396a# => X"b389c900",
		16#396b# => X"63e89d00",
		16#396c# => X"13840600",
		16#396d# => X"63949d04",
		16#396e# => X"63723c05",
		16#396f# => X"330cac01",
		16#3970# => X"3337ac01",
		16#3971# => X"33079701",
		16#3972# => X"b38ded00",
		16#3973# => X"1384f6ff",
		16#3974# => X"63e6bc01",
		16#3975# => X"6394bc03",
		16#3976# => X"6362ac03",
		16#3977# => X"63e69d00",
		16#3978# => X"639eb401",
		16#3979# => X"637c3c01",
		16#397a# => X"330cac01",
		16#397b# => X"3337ac01",
		16#397c# => X"33079701",
		16#397d# => X"1384e6ff",
		16#397e# => X"b38ded00",
		16#397f# => X"b3093c41",
		16#3980# => X"b3849d40",
		16#3981# => X"b3373c01",
		16#3982# => X"b384f440",
		16#3983# => X"9305f0ff",
		16#3984# => X"63889c1a",
		16#3985# => X"93850a00",
		16#3986# => X"13850400",
		16#3987# => X"ef400004",
		16#3988# => X"93050500",
		16#3989# => X"2324a100",
		16#398a# => X"13950c01",
		16#398b# => X"13550501",
		16#398c# => X"ef400000",
		16#398d# => X"2322a100",
		16#398e# => X"93850a00",
		16#398f# => X"13850400",
		16#3990# => X"ef404006",
		16#3991# => X"83268100",
		16#3992# => X"03274100",
		16#3993# => X"13150501",
		16#3994# => X"93d70901",
		16#3995# => X"33e5a700",
		16#3996# => X"938d0600",
		16#3997# => X"637ee500",
		16#3998# => X"33059501",
		16#3999# => X"938df6ff",
		16#399a# => X"63689501",
		16#399b# => X"6376e500",
		16#399c# => X"938de6ff",
		16#399d# => X"33059501",
		16#399e# => X"b304e540",
		16#399f# => X"93850a00",
		16#39a0# => X"13850400",
		16#39a1# => X"ef30907d",
		16#39a2# => X"93050500",
		16#39a3# => X"2322a100",
		16#39a4# => X"13950c01",
		16#39a5# => X"13550501",
		16#39a6# => X"ef309079",
		16#39a7# => X"130c0500",
		16#39a8# => X"93850a00",
		16#39a9# => X"13850400",
		16#39aa# => X"ef30d07f",
		16#39ab# => X"93990901",
		16#39ac# => X"03274100",
		16#39ad# => X"13150501",
		16#39ae# => X"93d90901",
		16#39af# => X"33e5a900",
		16#39b0# => X"93070700",
		16#39b1# => X"637e8501",
		16#39b2# => X"33059501",
		16#39b3# => X"9307f7ff",
		16#39b4# => X"63689501",
		16#39b5# => X"63768501",
		16#39b6# => X"9307e7ff",
		16#39b7# => X"33059501",
		16#39b8# => X"93940d01",
		16#39b9# => X"b3e4f400",
		16#39ba# => X"93970401",
		16#39bb# => X"93d70701",
		16#39bc# => X"93050b00",
		16#39bd# => X"b3098541",
		16#39be# => X"13850700",
		16#39bf# => X"2322f100",
		16#39c0# => X"93dd0401",
		16#39c1# => X"ef30d072",
		16#39c2# => X"93050b00",
		16#39c3# => X"930a0500",
		16#39c4# => X"13850d00",
		16#39c5# => X"ef30d071",
		16#39c6# => X"130c0500",
		16#39c7# => X"93850d00",
		16#39c8# => X"13850b00",
		16#39c9# => X"ef30d070",
		16#39ca# => X"83274100",
		16#39cb# => X"130b0500",
		16#39cc# => X"13850b00",
		16#39cd# => X"93850700",
		16#39ce# => X"ef30906f",
		16#39cf# => X"33058501",
		16#39d0# => X"93d70a01",
		16#39d1# => X"3385a700",
		16#39d2# => X"63768501",
		16#39d3# => X"b7070100",
		16#39d4# => X"330bfb00",
		16#39d5# => X"b7060100",
		16#39d6# => X"9386f6ff",
		16#39d7# => X"93570501",
		16#39d8# => X"3377d500",
		16#39d9# => X"13170701",
		16#39da# => X"b3fada00",
		16#39db# => X"b3876701",
		16#39dc# => X"33075701",
		16#39dd# => X"63e8f900",
		16#39de# => X"93850400",
		16#39df# => X"6390f904",
		16#39e0# => X"63000704",
		16#39e1# => X"33853c01",
		16#39e2# => X"9385f4ff",
		16#39e3# => X"63649503",
		16#39e4# => X"6366f500",
		16#39e5# => X"6314f502",
		16#39e6# => X"6370ed02",
		16#39e7# => X"93161d00",
		16#39e8# => X"33bda601",
		16#39e9# => X"b30c9d01",
		16#39ea# => X"9385e4ff",
		16#39eb# => X"33059501",
		16#39ec# => X"138d0600",
		16#39ed# => X"6314f500",
		16#39ee# => X"6304a701",
		16#39ef# => X"93e51500",
		16#39f0# => X"1307fa3f",
		16#39f1# => X"6352e012",
		16#39f2# => X"93f77500",
		16#39f3# => X"63800702",
		16#39f4# => X"93f7f500",
		16#39f5# => X"93064000",
		16#39f6# => X"638ad700",
		16#39f7# => X"93864500",
		16#39f8# => X"b3b5b600",
		16#39f9# => X"3304b400",
		16#39fa# => X"93850600",
		16#39fb# => X"93177400",
		16#39fc# => X"63da0700",
		16#39fd# => X"b70700ff",
		16#39fe# => X"9387f7ff",
		16#39ff# => X"3374f400",
		16#3a00# => X"13070a40",
		16#3a01# => X"9307e07f",
		16#3a02# => X"63c2e71a",
		16#3a03# => X"9317d401",
		16#3a04# => X"93d53500",
		16#3a05# => X"b3e7b700",
		16#3a06# => X"13543400",
		16#3a07# => X"b7061000",
		16#3a08# => X"9386f6ff",
		16#3a09# => X"3374d400",
		16#3a0a# => X"b7061080",
		16#3a0b# => X"1377f77f",
		16#3a0c# => X"9386f6ff",
		16#3a0d# => X"13174701",
		16#3a0e# => X"3374d400",
		16#3a0f# => X"1319f901",
		16#3a10# => X"3364e400",
		16#3a11# => X"33672401",
		16#3a12# => X"8320c104",
		16#3a13# => X"03248104",
		16#3a14# => X"83244104",
		16#3a15# => X"03290104",
		16#3a16# => X"8329c103",
		16#3a17# => X"032a8103",
		16#3a18# => X"832a4103",
		16#3a19# => X"032b0103",
		16#3a1a# => X"832bc102",
		16#3a1b# => X"032c8102",
		16#3a1c# => X"832c4102",
		16#3a1d# => X"032d0102",
		16#3a1e# => X"832dc101",
		16#3a1f# => X"13850700",
		16#3a20# => X"93050700",
		16#3a21# => X"13010105",
		16#3a22# => X"67800000",
		16#3a23# => X"130afaff",
		16#3a24# => X"130c0000",
		16#3a25# => X"6ff01fb9",
		16#3a26# => X"13890900",
		16#3a27# => X"13040b00",
		16#3a28# => X"93850400",
		16#3a29# => X"93870b00",
		16#3a2a# => X"13072000",
		16#3a2b# => X"6380e710",
		16#3a2c# => X"13073000",
		16#3a2d# => X"6382e70e",
		16#3a2e# => X"13071000",
		16#3a2f# => X"e392e7f0",
		16#3a30# => X"13040000",
		16#3a31# => X"93070000",
		16#3a32# => X"6f004009",
		16#3a33# => X"13890a00",
		16#3a34# => X"6ff09ffd",
		16#3a35# => X"37040800",
		16#3a36# => X"93050000",
		16#3a37# => X"13090000",
		16#3a38# => X"93073000",
		16#3a39# => X"6ff05ffc",
		16#3a3a# => X"93061000",
		16#3a3b# => X"b386e640",
		16#3a3c# => X"93078003",
		16#3a3d# => X"e3c6d7fc",
		16#3a3e# => X"9307f001",
		16#3a3f# => X"63c4d706",
		16#3a40# => X"130aea41",
		16#3a41# => X"b3174401",
		16#3a42# => X"33d7d500",
		16#3a43# => X"339a4501",
		16#3a44# => X"b3e7e700",
		16#3a45# => X"333a4001",
		16#3a46# => X"b3e74701",
		16#3a47# => X"3354d400",
		16#3a48# => X"13f77700",
		16#3a49# => X"63000702",
		16#3a4a# => X"13f7f700",
		16#3a4b# => X"93064000",
		16#3a4c# => X"630ad700",
		16#3a4d# => X"13874700",
		16#3a4e# => X"b337f700",
		16#3a4f# => X"3304f400",
		16#3a50# => X"93070700",
		16#3a51# => X"13178400",
		16#3a52# => X"634a0706",
		16#3a53# => X"1317d401",
		16#3a54# => X"93d73700",
		16#3a55# => X"b367f700",
		16#3a56# => X"13543400",
		16#3a57# => X"13070000",
		16#3a58# => X"6ff0dfeb",
		16#3a59# => X"930710fe",
		16#3a5a# => X"b387e740",
		16#3a5b# => X"13070002",
		16#3a5c# => X"b357f400",
		16#3a5d# => X"13050000",
		16#3a5e# => X"6386e600",
		16#3a5f# => X"130aea43",
		16#3a60# => X"33154401",
		16#3a61# => X"336ab500",
		16#3a62# => X"333a4001",
		16#3a63# => X"b3e74701",
		16#3a64# => X"13040000",
		16#3a65# => X"6ff0dff8",
		16#3a66# => X"37040800",
		16#3a67# => X"93070000",
		16#3a68# => X"1307f07f",
		16#3a69# => X"13090000",
		16#3a6a# => X"6ff05fe7",
		16#3a6b# => X"13040000",
		16#3a6c# => X"93070000",
		16#3a6d# => X"1307f07f",
		16#3a6e# => X"6ff05fe6",
		16#3a6f# => X"13040000",
		16#3a70# => X"93070000",
		16#3a71# => X"13071000",
		16#3a72# => X"6ff05fe5",
		16#3a73# => X"130101fa",
		16#3a74# => X"232c8104",
		16#3a75# => X"23263105",
		16#3a76# => X"37041000",
		16#3a77# => X"93d94501",
		16#3a78# => X"232a9104",
		16#3a79# => X"23206105",
		16#3a7a# => X"232e7103",
		16#3a7b# => X"232c8103",
		16#3a7c# => X"1304f4ff",
		16#3a7d# => X"232e1104",
		16#3a7e# => X"23282105",
		16#3a7f# => X"23244105",
		16#3a80# => X"23225105",
		16#3a81# => X"232a9103",
		16#3a82# => X"2328a103",
		16#3a83# => X"2326b103",
		16#3a84# => X"93f9f97f",
		16#3a85# => X"93040500",
		16#3a86# => X"930b0600",
		16#3a87# => X"138c0600",
		16#3a88# => X"3374b400",
		16#3a89# => X"13dbf501",
		16#3a8a# => X"6386090a",
		16#3a8b# => X"9307f07f",
		16#3a8c# => X"6384f910",
		16#3a8d# => X"37098000",
		16#3a8e# => X"13143400",
		16#3a8f# => X"33642401",
		16#3a90# => X"1359d501",
		16#3a91# => X"33698900",
		16#3a92# => X"131d3500",
		16#3a93# => X"938919c0",
		16#3a94# => X"930c0000",
		16#3a95# => X"13554c01",
		16#3a96# => X"370a1000",
		16#3a97# => X"130afaff",
		16#3a98# => X"1375f57f",
		16#3a99# => X"337a8a01",
		16#3a9a# => X"93840b00",
		16#3a9b# => X"135cfc01",
		16#3a9c# => X"63020510",
		16#3a9d# => X"9307f07f",
		16#3a9e# => X"6302f516",
		16#3a9f# => X"37048000",
		16#3aa0# => X"131a3a00",
		16#3aa1# => X"336a8a00",
		16#3aa2# => X"13d4db01",
		16#3aa3# => X"33644401",
		16#3aa4# => X"93943b00",
		16#3aa5# => X"130515c0",
		16#3aa6# => X"93070000",
		16#3aa7# => X"13972c00",
		16#3aa8# => X"3367f700",
		16#3aa9# => X"b389a900",
		16#3aaa# => X"1307f7ff",
		16#3aab# => X"9306e000",
		16#3aac# => X"b34b8b01",
		16#3aad# => X"938a1900",
		16#3aae# => X"63eee614",
		16#3aaf# => X"b7460110",
		16#3ab0# => X"13172700",
		16#3ab1# => X"93864664",
		16#3ab2# => X"3307d700",
		16#3ab3# => X"03270700",
		16#3ab4# => X"67000700",
		16#3ab5# => X"3369a400",
		16#3ab6# => X"630e0906",
		16#3ab7# => X"63000404",
		16#3ab8# => X"13050400",
		16#3ab9# => X"ef305042",
		16#3aba# => X"930755ff",
		16#3abb# => X"1307c001",
		16#3abc# => X"634cf702",
		16#3abd# => X"1309d001",
		16#3abe# => X"130d85ff",
		16#3abf# => X"3309f940",
		16#3ac0# => X"3314a401",
		16#3ac1# => X"33d92401",
		16#3ac2# => X"33698900",
		16#3ac3# => X"339da401",
		16#3ac4# => X"9309d0c0",
		16#3ac5# => X"b389a940",
		16#3ac6# => X"6ff09ff3",
		16#3ac7# => X"ef30d03e",
		16#3ac8# => X"13050502",
		16#3ac9# => X"6ff05ffc",
		16#3aca# => X"130985fd",
		16#3acb# => X"33992401",
		16#3acc# => X"130d0000",
		16#3acd# => X"6ff0dffd",
		16#3ace# => X"3369a400",
		16#3acf# => X"63040902",
		16#3ad0# => X"130d0500",
		16#3ad1# => X"13090400",
		16#3ad2# => X"9309f07f",
		16#3ad3# => X"930c3000",
		16#3ad4# => X"6ff05ff0",
		16#3ad5# => X"130d0000",
		16#3ad6# => X"93090000",
		16#3ad7# => X"930c1000",
		16#3ad8# => X"6ff05fef",
		16#3ad9# => X"130d0000",
		16#3ada# => X"9309f07f",
		16#3adb# => X"930c2000",
		16#3adc# => X"6ff05fee",
		16#3add# => X"33647a01",
		16#3ade# => X"630e0406",
		16#3adf# => X"63000a04",
		16#3ae0# => X"13050a00",
		16#3ae1# => X"ef305038",
		16#3ae2# => X"930755ff",
		16#3ae3# => X"1307c001",
		16#3ae4# => X"634ef702",
		16#3ae5# => X"1304d001",
		16#3ae6# => X"930485ff",
		16#3ae7# => X"3304f440",
		16#3ae8# => X"331a9a00",
		16#3ae9# => X"33d48b00",
		16#3aea# => X"33644401",
		16#3aeb# => X"b3949b00",
		16#3aec# => X"9307d0c0",
		16#3aed# => X"3385a740",
		16#3aee# => X"6ff01fee",
		16#3aef# => X"13850b00",
		16#3af0# => X"ef309034",
		16#3af1# => X"13050502",
		16#3af2# => X"6ff01ffc",
		16#3af3# => X"130485fd",
		16#3af4# => X"33948b00",
		16#3af5# => X"93040000",
		16#3af6# => X"6ff09ffd",
		16#3af7# => X"33647a01",
		16#3af8# => X"63020402",
		16#3af9# => X"13040a00",
		16#3afa# => X"1305f07f",
		16#3afb# => X"93073000",
		16#3afc# => X"6ff0dfea",
		16#3afd# => X"93040000",
		16#3afe# => X"13050000",
		16#3aff# => X"93071000",
		16#3b00# => X"6ff0dfe9",
		16#3b01# => X"93040000",
		16#3b02# => X"1305f07f",
		16#3b03# => X"93072000",
		16#3b04# => X"6ff0dfe8",
		16#3b05# => X"37070100",
		16#3b06# => X"130af7ff",
		16#3b07# => X"135c0d01",
		16#3b08# => X"93dd0401",
		16#3b09# => X"337d4d01",
		16#3b0a# => X"b3f44401",
		16#3b0b# => X"93050d00",
		16#3b0c# => X"13850400",
		16#3b0d# => X"2328e100",
		16#3b0e# => X"ef30901f",
		16#3b0f# => X"930c0500",
		16#3b10# => X"93850400",
		16#3b11# => X"13050c00",
		16#3b12# => X"ef30901e",
		16#3b13# => X"2326a100",
		16#3b14# => X"93850d00",
		16#3b15# => X"13050c00",
		16#3b16# => X"ef30901d",
		16#3b17# => X"130b0500",
		16#3b18# => X"93050d00",
		16#3b19# => X"13850d00",
		16#3b1a# => X"ef30901c",
		16#3b1b# => X"8326c100",
		16#3b1c# => X"93d70c01",
		16#3b1d# => X"3305d500",
		16#3b1e# => X"3385a700",
		16#3b1f# => X"6376d500",
		16#3b20# => X"03270101",
		16#3b21# => X"330beb00",
		16#3b22# => X"93560501",
		16#3b23# => X"33754501",
		16#3b24# => X"b3fc4c01",
		16#3b25# => X"13150501",
		16#3b26# => X"b3079501",
		16#3b27# => X"935c0401",
		16#3b28# => X"33744401",
		16#3b29# => X"93050d00",
		16#3b2a# => X"13050400",
		16#3b2b# => X"232ad100",
		16#3b2c# => X"2326f100",
		16#3b2d# => X"ef30d017",
		16#3b2e# => X"2328a100",
		16#3b2f# => X"93050400",
		16#3b30# => X"13050c00",
		16#3b31# => X"ef30d016",
		16#3b32# => X"130a0500",
		16#3b33# => X"93850c00",
		16#3b34# => X"13050c00",
		16#3b35# => X"ef30d015",
		16#3b36# => X"130c0500",
		16#3b37# => X"93050d00",
		16#3b38# => X"13850c00",
		16#3b39# => X"ef30d014",
		16#3b3a# => X"03270101",
		16#3b3b# => X"33054501",
		16#3b3c# => X"83264101",
		16#3b3d# => X"93570701",
		16#3b3e# => X"3385a700",
		16#3b3f# => X"63764501",
		16#3b40# => X"b7070100",
		16#3b41# => X"330cfc00",
		16#3b42# => X"37060100",
		16#3b43# => X"93570501",
		16#3b44# => X"338c8701",
		16#3b45# => X"9307f6ff",
		16#3b46# => X"337af500",
		16#3b47# => X"3377f700",
		16#3b48# => X"131a0a01",
		16#3b49# => X"135d0901",
		16#3b4a# => X"330aea00",
		16#3b4b# => X"3379f900",
		16#3b4c# => X"33874601",
		16#3b4d# => X"93050900",
		16#3b4e# => X"13850400",
		16#3b4f# => X"2328e100",
		16#3b50# => X"232ec100",
		16#3b51# => X"ef30d00e",
		16#3b52# => X"93850400",
		16#3b53# => X"232ca100",
		16#3b54# => X"13050d00",
		16#3b55# => X"ef30d00d",
		16#3b56# => X"232aa100",
		16#3b57# => X"93050d00",
		16#3b58# => X"13850d00",
		16#3b59# => X"ef30d00c",
		16#3b5a# => X"93040500",
		16#3b5b# => X"93050900",
		16#3b5c# => X"13850d00",
		16#3b5d# => X"ef30d00b",
		16#3b5e# => X"83264101",
		16#3b5f# => X"03278101",
		16#3b60# => X"3305d500",
		16#3b61# => X"93570701",
		16#3b62# => X"3385a700",
		16#3b63# => X"6376d500",
		16#3b64# => X"0326c101",
		16#3b65# => X"b384c400",
		16#3b66# => X"b7060100",
		16#3b67# => X"9387f6ff",
		16#3b68# => X"935d0501",
		16#3b69# => X"b3849d00",
		16#3b6a# => X"b37df500",
		16#3b6b# => X"3377f700",
		16#3b6c# => X"93050900",
		16#3b6d# => X"13050400",
		16#3b6e# => X"939d0d01",
		16#3b6f# => X"b38ded00",
		16#3b70# => X"232cd100",
		16#3b71# => X"ef30d006",
		16#3b72# => X"93050400",
		16#3b73# => X"232aa100",
		16#3b74# => X"13050d00",
		16#3b75# => X"ef30d005",
		16#3b76# => X"93050d00",
		16#3b77# => X"13040500",
		16#3b78# => X"13850c00",
		16#3b79# => X"ef30d004",
		16#3b7a# => X"130d0500",
		16#3b7b# => X"93050900",
		16#3b7c# => X"13850c00",
		16#3b7d# => X"ef30d003",
		16#3b7e# => X"03274101",
		16#3b7f# => X"33058500",
		16#3b80# => X"93570701",
		16#3b81# => X"3385a700",
		16#3b82# => X"63768500",
		16#3b83# => X"83268101",
		16#3b84# => X"330ddd00",
		16#3b85# => X"83270101",
		16#3b86# => X"b7060100",
		16#3b87# => X"9386f6ff",
		16#3b88# => X"330bfb00",
		16#3b89# => X"b377d500",
		16#3b8a# => X"3377d700",
		16#3b8b# => X"93970701",
		16#3b8c# => X"b387e700",
		16#3b8d# => X"333a4b01",
		16#3b8e# => X"b3878701",
		16#3b8f# => X"33844701",
		16#3b90# => X"330bbb01",
		16#3b91# => X"33079400",
		16#3b92# => X"b33dbb01",
		16#3b93# => X"b306b701",
		16#3b94# => X"33bc8701",
		16#3b95# => X"33344401",
		16#3b96# => X"93570501",
		16#3b97# => X"33379700",
		16#3b98# => X"33648c00",
		16#3b99# => X"b3bdb601",
		16#3b9a# => X"3304f400",
		16#3b9b# => X"b36db701",
		16#3b9c# => X"3304b401",
		16#3b9d# => X"3304a401",
		16#3b9e# => X"93d77601",
		16#3b9f# => X"13149400",
		16#3ba0# => X"3364f400",
		16#3ba1# => X"8327c100",
		16#3ba2# => X"93149b00",
		16#3ba3# => X"135b7b01",
		16#3ba4# => X"b3e4f400",
		16#3ba5# => X"b3349000",
		16#3ba6# => X"93979600",
		16#3ba7# => X"b3e46401",
		16#3ba8# => X"b3e4f400",
		16#3ba9# => X"93177400",
		16#3baa# => X"63d20712",
		16#3bab# => X"93d71400",
		16#3bac# => X"93f41400",
		16#3bad# => X"b3e49700",
		16#3bae# => X"9317f401",
		16#3baf# => X"b3e4f400",
		16#3bb0# => X"13541400",
		16#3bb1# => X"1387fa3f",
		16#3bb2# => X"6356e010",
		16#3bb3# => X"93f77400",
		16#3bb4# => X"63800702",
		16#3bb5# => X"93f7f400",
		16#3bb6# => X"93064000",
		16#3bb7# => X"638ad700",
		16#3bb8# => X"93874400",
		16#3bb9# => X"b3b49700",
		16#3bba# => X"33049400",
		16#3bbb# => X"93840700",
		16#3bbc# => X"93177400",
		16#3bbd# => X"63da0700",
		16#3bbe# => X"b70700ff",
		16#3bbf# => X"9387f7ff",
		16#3bc0# => X"3374f400",
		16#3bc1# => X"13870a40",
		16#3bc2# => X"9307e07f",
		16#3bc3# => X"63c6e718",
		16#3bc4# => X"93da3400",
		16#3bc5# => X"9314d401",
		16#3bc6# => X"b3e45401",
		16#3bc7# => X"13543400",
		16#3bc8# => X"b7071000",
		16#3bc9# => X"9387f7ff",
		16#3bca# => X"3374f400",
		16#3bcb# => X"9377f77f",
		16#3bcc# => X"37071080",
		16#3bcd# => X"1307f7ff",
		16#3bce# => X"93974701",
		16#3bcf# => X"3374e400",
		16#3bd0# => X"939bfb01",
		16#3bd1# => X"3364f400",
		16#3bd2# => X"b3677401",
		16#3bd3# => X"8320c105",
		16#3bd4# => X"03248105",
		16#3bd5# => X"13850400",
		16#3bd6# => X"03290105",
		16#3bd7# => X"83244105",
		16#3bd8# => X"8329c104",
		16#3bd9# => X"032a8104",
		16#3bda# => X"832a4104",
		16#3bdb# => X"032b0104",
		16#3bdc# => X"832bc103",
		16#3bdd# => X"032c8103",
		16#3bde# => X"832c4103",
		16#3bdf# => X"032d0103",
		16#3be0# => X"832dc102",
		16#3be1# => X"93850700",
		16#3be2# => X"13010106",
		16#3be3# => X"67800000",
		16#3be4# => X"930b0b00",
		16#3be5# => X"13040900",
		16#3be6# => X"93040d00",
		16#3be7# => X"93870c00",
		16#3be8# => X"13072000",
		16#3be9# => X"638ae70e",
		16#3bea# => X"13073000",
		16#3beb# => X"638ce70c",
		16#3bec# => X"13071000",
		16#3bed# => X"e398e7f0",
		16#3bee# => X"13040000",
		16#3bef# => X"93040000",
		16#3bf0# => X"6f008008",
		16#3bf1# => X"930b0c00",
		16#3bf2# => X"6ff09ffd",
		16#3bf3# => X"938a0900",
		16#3bf4# => X"6ff05fef",
		16#3bf5# => X"93061000",
		16#3bf6# => X"b386e640",
		16#3bf7# => X"93078003",
		16#3bf8# => X"e3ccd7fc",
		16#3bf9# => X"9307f001",
		16#3bfa# => X"63c4d706",
		16#3bfb# => X"938aea41",
		16#3bfc# => X"b3175401",
		16#3bfd# => X"33d7d400",
		16#3bfe# => X"b3945401",
		16#3bff# => X"b3e7e700",
		16#3c00# => X"b3349000",
		16#3c01# => X"b3e49700",
		16#3c02# => X"3354d400",
		16#3c03# => X"93f77400",
		16#3c04# => X"63800702",
		16#3c05# => X"93f7f400",
		16#3c06# => X"13074000",
		16#3c07# => X"638ae700",
		16#3c08# => X"93874400",
		16#3c09# => X"b3b49700",
		16#3c0a# => X"33049400",
		16#3c0b# => X"93840700",
		16#3c0c# => X"93178400",
		16#3c0d# => X"63ca0706",
		16#3c0e# => X"9317d401",
		16#3c0f# => X"93d43400",
		16#3c10# => X"b3e49700",
		16#3c11# => X"13543400",
		16#3c12# => X"13070000",
		16#3c13# => X"6ff05fed",
		16#3c14# => X"930710fe",
		16#3c15# => X"b387e740",
		16#3c16# => X"13060002",
		16#3c17# => X"b357f400",
		16#3c18# => X"13070000",
		16#3c19# => X"6386c600",
		16#3c1a# => X"938aea43",
		16#3c1b# => X"33175401",
		16#3c1c# => X"b3649700",
		16#3c1d# => X"b3349000",
		16#3c1e# => X"b3e49700",
		16#3c1f# => X"13040000",
		16#3c20# => X"6ff0dff8",
		16#3c21# => X"37040800",
		16#3c22# => X"93040000",
		16#3c23# => X"1307f07f",
		16#3c24# => X"930b0000",
		16#3c25# => X"6ff0dfe8",
		16#3c26# => X"13040000",
		16#3c27# => X"93040000",
		16#3c28# => X"1307f07f",
		16#3c29# => X"6ff0dfe7",
		16#3c2a# => X"13040000",
		16#3c2b# => X"93040000",
		16#3c2c# => X"13071000",
		16#3c2d# => X"6ff0dfe6",
		16#3c2e# => X"8327c500",
		16#3c2f# => X"03af0500",
		16#3c30# => X"83af4500",
		16#3c31# => X"83a28500",
		16#3c32# => X"83a5c500",
		16#3c33# => X"37870000",
		16#3c34# => X"93d60701",
		16#3c35# => X"1307f7ff",
		16#3c36# => X"13980701",
		16#3c37# => X"939e0501",
		16#3c38# => X"13d6f701",
		16#3c39# => X"b3f6e600",
		16#3c3a# => X"93d70501",
		16#3c3b# => X"130101ff",
		16#3c3c# => X"83280500",
		16#3c3d# => X"03234500",
		16#3c3e# => X"032e8500",
		16#3c3f# => X"13580801",
		16#3c40# => X"93de0e01",
		16#3c41# => X"b3f7e700",
		16#3c42# => X"93d5f501",
		16#3c43# => X"6390e602",
		16#3c44# => X"33e76800",
		16#3c45# => X"3367c701",
		16#3c46# => X"33670701",
		16#3c47# => X"13051000",
		16#3c48# => X"631a0704",
		16#3c49# => X"6398d704",
		16#3c4a# => X"6f008000",
		16#3c4b# => X"639ce700",
		16#3c4c# => X"3367ff01",
		16#3c4d# => X"33675700",
		16#3c4e# => X"3367d701",
		16#3c4f# => X"13051000",
		16#3c50# => X"631a0702",
		16#3c51# => X"13051000",
		16#3c52# => X"6396d702",
		16#3c53# => X"6394e803",
		16#3c54# => X"6312f303",
		16#3c55# => X"63105e02",
		16#3c56# => X"631ed801",
		16#3c57# => X"6300b602",
		16#3c58# => X"639a0700",
		16#3c59# => X"33e56800",
		16#3c5a# => X"3365c501",
		16#3c5b# => X"33650501",
		16#3c5c# => X"3335a000",
		16#3c5d# => X"13010101",
		16#3c5e# => X"67800000",
		16#3c5f# => X"13050000",
		16#3c60# => X"6ff05fff",
		16#3c61# => X"8327c500",
		16#3c62# => X"83a8c500",
		16#3c63# => X"032f0500",
		16#3c64# => X"03264500",
		16#3c65# => X"03288500",
		16#3c66# => X"37850000",
		16#3c67# => X"13d70701",
		16#3c68# => X"1305f5ff",
		16#3c69# => X"939e0801",
		16#3c6a# => X"93d60801",
		16#3c6b# => X"83a20500",
		16#3c6c# => X"03a34500",
		16#3c6d# => X"03ae8500",
		16#3c6e# => X"3377a700",
		16#3c6f# => X"93950701",
		16#3c70# => X"130101ff",
		16#3c71# => X"93d50501",
		16#3c72# => X"93d7f701",
		16#3c73# => X"93de0e01",
		16#3c74# => X"b3f6a600",
		16#3c75# => X"93d8f801",
		16#3c76# => X"6310a702",
		16#3c77# => X"b36fcf00",
		16#3c78# => X"b3ef0f01",
		16#3c79# => X"b3efbf00",
		16#3c7a# => X"1305e0ff",
		16#3c7b# => X"63800f0e",
		16#3c7c# => X"13010101",
		16#3c7d# => X"67800000",
		16#3c7e# => X"6398a602",
		16#3c7f# => X"b3ef6200",
		16#3c80# => X"b3efcf01",
		16#3c81# => X"b3efdf01",
		16#3c82# => X"1305e0ff",
		16#3c83# => X"e3920ffe",
		16#3c84# => X"63120704",
		16#3c85# => X"3365cf00",
		16#3c86# => X"33650501",
		16#3c87# => X"3365b500",
		16#3c88# => X"13351500",
		16#3c89# => X"6f00c002",
		16#3c8a# => X"6314070a",
		16#3c8b# => X"3365cf00",
		16#3c8c# => X"33650501",
		16#3c8d# => X"3365b500",
		16#3c8e# => X"13351500",
		16#3c8f# => X"639a0600",
		16#3c90# => X"b3ef6200",
		16#3c91# => X"b3efcf01",
		16#3c92# => X"b3efdf01",
		16#3c93# => X"638c0f06",
		16#3c94# => X"631a0500",
		16#3c95# => X"638e1701",
		16#3c96# => X"13051000",
		16#3c97# => X"e38a07f8",
		16#3c98# => X"6f008000",
		16#3c99# => X"e39608f8",
		16#3c9a# => X"1305f0ff",
		16#3c9b# => X"6ff05ff8",
		16#3c9c# => X"e3c4e6fe",
		16#3c9d# => X"635ad700",
		16#3c9e# => X"1305f0ff",
		16#3c9f# => X"e38a07f6",
		16#3ca0# => X"13051000",
		16#3ca1# => X"6ff0dff6",
		16#3ca2# => X"e3e8befc",
		16#3ca3# => X"6396d503",
		16#3ca4# => X"e3640efd",
		16#3ca5# => X"6314c805",
		16#3ca6# => X"e360c3fc",
		16#3ca7# => X"63146600",
		16#3ca8# => X"e3ece2fb",
		16#3ca9# => X"e36a66fc",
		16#3caa# => X"13050000",
		16#3cab# => X"e31266f4",
		16#3cac# => X"e3645ffc",
		16#3cad# => X"6ff0dff3",
		16#3cae# => X"e3e0d5fd",
		16#3caf# => X"13050000",
		16#3cb0# => X"6ff01ff3",
		16#3cb1# => X"e31c05fe",
		16#3cb2# => X"6ff01ff9",
		16#3cb3# => X"e388e6f2",
		16#3cb4# => X"13050000",
		16#3cb5# => X"e38606f6",
		16#3cb6# => X"6ff0dff7",
		16#3cb7# => X"e36ec8f9",
		16#3cb8# => X"6ff0dffd",
		16#3cb9# => X"8327c500",
		16#3cba# => X"83a8c500",
		16#3cbb# => X"032f0500",
		16#3cbc# => X"03264500",
		16#3cbd# => X"03288500",
		16#3cbe# => X"37850000",
		16#3cbf# => X"13d70701",
		16#3cc0# => X"1305f5ff",
		16#3cc1# => X"939e0801",
		16#3cc2# => X"93d60801",
		16#3cc3# => X"83a20500",
		16#3cc4# => X"03a34500",
		16#3cc5# => X"03ae8500",
		16#3cc6# => X"3377a700",
		16#3cc7# => X"93950701",
		16#3cc8# => X"130101ff",
		16#3cc9# => X"93d50501",
		16#3cca# => X"93d7f701",
		16#3ccb# => X"93de0e01",
		16#3ccc# => X"b3f6a600",
		16#3ccd# => X"93d8f801",
		16#3cce# => X"6310a702",
		16#3ccf# => X"b36fcf00",
		16#3cd0# => X"b3ef0f01",
		16#3cd1# => X"b3efbf00",
		16#3cd2# => X"13052000",
		16#3cd3# => X"63800f0e",
		16#3cd4# => X"13010101",
		16#3cd5# => X"67800000",
		16#3cd6# => X"6398a602",
		16#3cd7# => X"b3ef6200",
		16#3cd8# => X"b3efcf01",
		16#3cd9# => X"b3efdf01",
		16#3cda# => X"13052000",
		16#3cdb# => X"e3920ffe",
		16#3cdc# => X"63120704",
		16#3cdd# => X"3365cf00",
		16#3cde# => X"33650501",
		16#3cdf# => X"3365b500",
		16#3ce0# => X"13351500",
		16#3ce1# => X"6f00c002",
		16#3ce2# => X"6314070a",
		16#3ce3# => X"3365cf00",
		16#3ce4# => X"33650501",
		16#3ce5# => X"3365b500",
		16#3ce6# => X"13351500",
		16#3ce7# => X"639a0600",
		16#3ce8# => X"b3ef6200",
		16#3ce9# => X"b3efcf01",
		16#3cea# => X"b3efdf01",
		16#3ceb# => X"638c0f06",
		16#3cec# => X"631a0500",
		16#3ced# => X"638e1701",
		16#3cee# => X"13051000",
		16#3cef# => X"e38a07f8",
		16#3cf0# => X"6f008000",
		16#3cf1# => X"e39608f8",
		16#3cf2# => X"1305f0ff",
		16#3cf3# => X"6ff05ff8",
		16#3cf4# => X"e3c4e6fe",
		16#3cf5# => X"635ad700",
		16#3cf6# => X"1305f0ff",
		16#3cf7# => X"e38a07f6",
		16#3cf8# => X"13051000",
		16#3cf9# => X"6ff0dff6",
		16#3cfa# => X"e3e8befc",
		16#3cfb# => X"6396d503",
		16#3cfc# => X"e3640efd",
		16#3cfd# => X"6314c805",
		16#3cfe# => X"e360c3fc",
		16#3cff# => X"63146600",
		16#3d00# => X"e3ece2fb",
		16#3d01# => X"e36a66fc",
		16#3d02# => X"13050000",
		16#3d03# => X"e31266f4",
		16#3d04# => X"e3645ffc",
		16#3d05# => X"6ff0dff3",
		16#3d06# => X"e3e0d5fd",
		16#3d07# => X"13050000",
		16#3d08# => X"6ff01ff3",
		16#3d09# => X"e31c05fe",
		16#3d0a# => X"6ff01ff9",
		16#3d0b# => X"e388e6f2",
		16#3d0c# => X"13050000",
		16#3d0d# => X"e38606f6",
		16#3d0e# => X"6ff0dff7",
		16#3d0f# => X"e36ec8f9",
		16#3d10# => X"6ff0dffd",
		16#3d11# => X"130101f2",
		16#3d12# => X"2326310d",
		16#3d13# => X"83a9c500",
		16#3d14# => X"83a60500",
		16#3d15# => X"83a74500",
		16#3d16# => X"2328a100",
		16#3d17# => X"03a58500",
		16#3d18# => X"13970901",
		16#3d19# => X"2328210d",
		16#3d1a# => X"2324410d",
		16#3d1b# => X"2322510d",
		16#3d1c# => X"2320610d",
		16#3d1d# => X"032a0600",
		16#3d1e# => X"032b4600",
		16#3d1f# => X"832a8600",
		16#3d20# => X"0329c600",
		16#3d21# => X"37860000",
		16#3d22# => X"232c810c",
		16#3d23# => X"13570701",
		16#3d24# => X"13d40901",
		16#3d25# => X"1306f6ff",
		16#3d26# => X"23263109",
		16#3d27# => X"232e110c",
		16#3d28# => X"232a910c",
		16#3d29# => X"232e710b",
		16#3d2a# => X"232c810b",
		16#3d2b# => X"232a910b",
		16#3d2c# => X"2328a10b",
		16#3d2d# => X"2326b10b",
		16#3d2e# => X"2320d108",
		16#3d2f# => X"2322f108",
		16#3d30# => X"2324a108",
		16#3d31# => X"2328d104",
		16#3d32# => X"232af104",
		16#3d33# => X"232ca104",
		16#3d34# => X"232ee104",
		16#3d35# => X"3374c400",
		16#3d36# => X"93d9f901",
		16#3d37# => X"63080412",
		16#3d38# => X"630ec424",
		16#3d39# => X"37050100",
		16#3d3a# => X"3365a700",
		16#3d3b# => X"232ea104",
		16#3d3c# => X"13060105",
		16#3d3d# => X"9307c105",
		16#3d3e# => X"03a70700",
		16#3d3f# => X"83a6c7ff",
		16#3d40# => X"9387c7ff",
		16#3d41# => X"13173700",
		16#3d42# => X"93d6d601",
		16#3d43# => X"3367d700",
		16#3d44# => X"23a2e700",
		16#3d45# => X"e312f6fe",
		16#3d46# => X"83270105",
		16#3d47# => X"93973700",
		16#3d48# => X"2328f104",
		16#3d49# => X"b7c7ffff",
		16#3d4a# => X"93871700",
		16#3d4b# => X"3304f400",
		16#3d4c# => X"93040000",
		16#3d4d# => X"93170901",
		16#3d4e# => X"37870000",
		16#3d4f# => X"13550901",
		16#3d50# => X"93d70701",
		16#3d51# => X"1307f7ff",
		16#3d52# => X"23262109",
		16#3d53# => X"23204109",
		16#3d54# => X"23226109",
		16#3d55# => X"23245109",
		16#3d56# => X"23204107",
		16#3d57# => X"23226107",
		16#3d58# => X"23245107",
		16#3d59# => X"2326f106",
		16#3d5a# => X"3375e500",
		16#3d5b# => X"1359f901",
		16#3d5c# => X"630a051e",
		16#3d5d# => X"6302e532",
		16#3d5e# => X"b70a0100",
		16#3d5f# => X"b3ea5701",
		16#3d60# => X"23265107",
		16#3d61# => X"13060106",
		16#3d62# => X"9307c106",
		16#3d63# => X"03a70700",
		16#3d64# => X"83a6c7ff",
		16#3d65# => X"9387c7ff",
		16#3d66# => X"13173700",
		16#3d67# => X"93d6d601",
		16#3d68# => X"3367d700",
		16#3d69# => X"23a2e700",
		16#3d6a# => X"e312f6fe",
		16#3d6b# => X"83270106",
		16#3d6c# => X"93973700",
		16#3d6d# => X"2320f106",
		16#3d6e# => X"b7c7ffff",
		16#3d6f# => X"93871700",
		16#3d70# => X"3305f500",
		16#3d71# => X"13070000",
		16#3d72# => X"b3c72901",
		16#3d73# => X"232af100",
		16#3d74# => X"b3078500",
		16#3d75# => X"2324f102",
		16#3d76# => X"93871700",
		16#3d77# => X"2322f102",
		16#3d78# => X"93972400",
		16#3d79# => X"b3e7e700",
		16#3d7a# => X"9387f7ff",
		16#3d7b# => X"9306e000",
		16#3d7c# => X"63e8f62c",
		16#3d7d# => X"b7460110",
		16#3d7e# => X"93972700",
		16#3d7f# => X"93860668",
		16#3d80# => X"b387d700",
		16#3d81# => X"83a70700",
		16#3d82# => X"67800700",
		16#3d83# => X"33e6d700",
		16#3d84# => X"3366a600",
		16#3d85# => X"3366e600",
		16#3d86# => X"63000614",
		16#3d87# => X"63020706",
		16#3d88# => X"13050700",
		16#3d89# => X"ef30400e",
		16#3d8a# => X"130c0500",
		16#3d8b# => X"930b4cff",
		16#3d8c# => X"93d45b40",
		16#3d8d# => X"93fbfb01",
		16#3d8e# => X"638e0b06",
		16#3d8f# => X"9305c0ff",
		16#3d90# => X"13850400",
		16#3d91# => X"ef20d07e",
		16#3d92# => X"93060002",
		16#3d93# => X"13972400",
		16#3d94# => X"130800ff",
		16#3d95# => X"b3867641",
		16#3d96# => X"1305c5ff",
		16#3d97# => X"63160509",
		16#3d98# => X"9307010a",
		16#3d99# => X"3387e700",
		16#3d9a# => X"83270105",
		16#3d9b# => X"9384f4ff",
		16#3d9c# => X"b39b7701",
		16#3d9d# => X"232877fb",
		16#3d9e# => X"1307f0ff",
		16#3d9f# => X"6f00c00a",
		16#3da0# => X"63080500",
		16#3da1# => X"ef304008",
		16#3da2# => X"130c0502",
		16#3da3# => X"6ff01ffa",
		16#3da4# => X"638a0700",
		16#3da5# => X"13850700",
		16#3da6# => X"ef300007",
		16#3da7# => X"130c0504",
		16#3da8# => X"6ff0dff8",
		16#3da9# => X"13850600",
		16#3daa# => X"ef300006",
		16#3dab# => X"130c0506",
		16#3dac# => X"6ff0dff7",
		16#3dad# => X"9305c0ff",
		16#3dae# => X"13850400",
		16#3daf# => X"ef205077",
		16#3db0# => X"13040105",
		16#3db1# => X"93073000",
		16#3db2# => X"3307a400",
		16#3db3# => X"0327c700",
		16#3db4# => X"9387f7ff",
		16#3db5# => X"1304c4ff",
		16#3db6# => X"2328e400",
		16#3db7# => X"e3d697fe",
		16#3db8# => X"9384f4ff",
		16#3db9# => X"6ff05ff9",
		16#3dba# => X"93070105",
		16#3dbb# => X"b385a700",
		16#3dbc# => X"3306a700",
		16#3dbd# => X"3386c700",
		16#3dbe# => X"83a7c500",
		16#3dbf# => X"83a50501",
		16#3dc0# => X"b3d7d700",
		16#3dc1# => X"b3957501",
		16#3dc2# => X"b3e7b700",
		16#3dc3# => X"2328f600",
		16#3dc4# => X"6ff09ff4",
		16#3dc5# => X"93972400",
		16#3dc6# => X"93060105",
		16#3dc7# => X"b387f600",
		16#3dc8# => X"23a00700",
		16#3dc9# => X"9384f4ff",
		16#3dca# => X"e396e4fe",
		16#3dcb# => X"37c4ffff",
		16#3dcc# => X"13041401",
		16#3dcd# => X"33048441",
		16#3dce# => X"6ff09fdf",
		16#3dcf# => X"b3e7d700",
		16#3dd0# => X"b3e7a700",
		16#3dd1# => X"33e5e700",
		16#3dd2# => X"93042000",
		16#3dd3# => X"e30405de",
		16#3dd4# => X"93043000",
		16#3dd5# => X"6ff01fde",
		16#3dd6# => X"13040000",
		16#3dd7# => X"93041000",
		16#3dd8# => X"6ff05fdd",
		16#3dd9# => X"33676a01",
		16#3dda# => X"33675701",
		16#3ddb# => X"3367f700",
		16#3ddc# => X"63020714",
		16#3ddd# => X"63820706",
		16#3dde# => X"13850700",
		16#3ddf# => X"ef20d078",
		16#3de0# => X"130b0500",
		16#3de1# => X"930a4bff",
		16#3de2# => X"13da5a40",
		16#3de3# => X"93fafa01",
		16#3de4# => X"63800a08",
		16#3de5# => X"9305c0ff",
		16#3de6# => X"13050a00",
		16#3de7# => X"ef205069",
		16#3de8# => X"93060002",
		16#3de9# => X"13172a00",
		16#3dea# => X"130800ff",
		16#3deb# => X"b3865641",
		16#3dec# => X"1305c5ff",
		16#3ded# => X"63180509",
		16#3dee# => X"9307010a",
		16#3def# => X"3387e700",
		16#3df0# => X"83270106",
		16#3df1# => X"130afaff",
		16#3df2# => X"b39a5701",
		16#3df3# => X"232057fd",
		16#3df4# => X"1307f0ff",
		16#3df5# => X"6f00000b",
		16#3df6# => X"638a0a00",
		16#3df7# => X"13850a00",
		16#3df8# => X"ef209072",
		16#3df9# => X"130b0502",
		16#3dfa# => X"6ff0dff9",
		16#3dfb# => X"630a0b00",
		16#3dfc# => X"13050b00",
		16#3dfd# => X"ef205071",
		16#3dfe# => X"130b0504",
		16#3dff# => X"6ff09ff8",
		16#3e00# => X"13050a00",
		16#3e01# => X"ef205070",
		16#3e02# => X"130b0506",
		16#3e03# => X"6ff09ff7",
		16#3e04# => X"9305c0ff",
		16#3e05# => X"13050a00",
		16#3e06# => X"ef209061",
		16#3e07# => X"930a0106",
		16#3e08# => X"93073000",
		16#3e09# => X"3387aa00",
		16#3e0a# => X"0327c700",
		16#3e0b# => X"9387f7ff",
		16#3e0c# => X"938acaff",
		16#3e0d# => X"23a8ea00",
		16#3e0e# => X"e3d647ff",
		16#3e0f# => X"130afaff",
		16#3e10# => X"6ff01ff9",
		16#3e11# => X"93070106",
		16#3e12# => X"b385a700",
		16#3e13# => X"3306a700",
		16#3e14# => X"3386c700",
		16#3e15# => X"83a7c500",
		16#3e16# => X"83a50501",
		16#3e17# => X"b3d7d700",
		16#3e18# => X"b3955501",
		16#3e19# => X"b3e7b700",
		16#3e1a# => X"2328f600",
		16#3e1b# => X"6ff05ff4",
		16#3e1c# => X"93172a00",
		16#3e1d# => X"93060106",
		16#3e1e# => X"b387f600",
		16#3e1f# => X"23a00700",
		16#3e20# => X"130afaff",
		16#3e21# => X"e316eafe",
		16#3e22# => X"37c5ffff",
		16#3e23# => X"13051501",
		16#3e24# => X"33056541",
		16#3e25# => X"6ff01fd3",
		16#3e26# => X"336a6a01",
		16#3e27# => X"b36a5a01",
		16#3e28# => X"b3eafa00",
		16#3e29# => X"13072000",
		16#3e2a# => X"e3800ad2",
		16#3e2b# => X"13073000",
		16#3e2c# => X"6ff09fd1",
		16#3e2d# => X"13050000",
		16#3e2e# => X"13071000",
		16#3e2f# => X"6ff0dfd0",
		16#3e30# => X"83290105",
		16#3e31# => X"03240106",
		16#3e32# => X"370b0100",
		16#3e33# => X"9304fbff",
		16#3e34# => X"93da0901",
		16#3e35# => X"13590401",
		16#3e36# => X"b3f99900",
		16#3e37# => X"33749400",
		16#3e38# => X"93850900",
		16#3e39# => X"13050400",
		16#3e3a# => X"ef209054",
		16#3e3b# => X"130a0500",
		16#3e3c# => X"93050400",
		16#3e3d# => X"13850a00",
		16#3e3e# => X"ef209053",
		16#3e3f# => X"130c0500",
		16#3e40# => X"93050900",
		16#3e41# => X"13850a00",
		16#3e42# => X"ef209052",
		16#3e43# => X"930b0500",
		16#3e44# => X"93850900",
		16#3e45# => X"13050900",
		16#3e46# => X"ef209051",
		16#3e47# => X"33058501",
		16#3e48# => X"93570a01",
		16#3e49# => X"3385a700",
		16#3e4a# => X"63748501",
		16#3e4b# => X"b38b6b01",
		16#3e4c# => X"832c4106",
		16#3e4d# => X"135d0501",
		16#3e4e# => X"33759500",
		16#3e4f# => X"337a9a00",
		16#3e50# => X"13150501",
		16#3e51# => X"b3074501",
		16#3e52# => X"13da0c01",
		16#3e53# => X"b3fc9c00",
		16#3e54# => X"93850900",
		16#3e55# => X"13850c00",
		16#3e56# => X"2326f102",
		16#3e57# => X"2320f108",
		16#3e58# => X"ef20104d",
		16#3e59# => X"130b0500",
		16#3e5a# => X"93850c00",
		16#3e5b# => X"13850a00",
		16#3e5c# => X"ef20104c",
		16#3e5d# => X"93040500",
		16#3e5e# => X"93050a00",
		16#3e5f# => X"13850a00",
		16#3e60# => X"ef20104b",
		16#3e61# => X"130c0500",
		16#3e62# => X"93850900",
		16#3e63# => X"13050a00",
		16#3e64# => X"ef20104a",
		16#3e65# => X"33059500",
		16#3e66# => X"93570b01",
		16#3e67# => X"3385a700",
		16#3e68# => X"63769500",
		16#3e69# => X"b7070100",
		16#3e6a# => X"330cfc00",
		16#3e6b# => X"b7060100",
		16#3e6c# => X"93570501",
		16#3e6d# => X"232cf100",
		16#3e6e# => X"9387f6ff",
		16#3e6f# => X"b37df500",
		16#3e70# => X"83244105",
		16#3e71# => X"337bfb00",
		16#3e72# => X"939d0d01",
		16#3e73# => X"b38d6d01",
		16#3e74# => X"3307bd01",
		16#3e75# => X"13dd0401",
		16#3e76# => X"b3f4f400",
		16#3e77# => X"93850400",
		16#3e78# => X"13050400",
		16#3e79# => X"232ae102",
		16#3e7a# => X"2324d100",
		16#3e7b# => X"ef205044",
		16#3e7c# => X"2322a100",
		16#3e7d# => X"93050400",
		16#3e7e# => X"13050d00",
		16#3e7f# => X"ef205043",
		16#3e80# => X"2320a100",
		16#3e81# => X"93050d00",
		16#3e82# => X"13050900",
		16#3e83# => X"ef205042",
		16#3e84# => X"130b0500",
		16#3e85# => X"93850400",
		16#3e86# => X"13050900",
		16#3e87# => X"ef205041",
		16#3e88# => X"03260100",
		16#3e89# => X"03274100",
		16#3e8a# => X"3305c500",
		16#3e8b# => X"93570701",
		16#3e8c# => X"3385a700",
		16#3e8d# => X"6376c500",
		16#3e8e# => X"83268100",
		16#3e8f# => X"330bdb00",
		16#3e90# => X"93570501",
		16#3e91# => X"37060100",
		16#3e92# => X"b3876701",
		16#3e93# => X"232ef100",
		16#3e94# => X"9307f6ff",
		16#3e95# => X"337bf500",
		16#3e96# => X"3377f700",
		16#3e97# => X"93850c00",
		16#3e98# => X"131b0b01",
		16#3e99# => X"13850400",
		16#3e9a# => X"330beb00",
		16#3e9b# => X"2326c100",
		16#3e9c# => X"ef20103c",
		16#3e9d# => X"2324a100",
		16#3e9e# => X"93850c00",
		16#3e9f# => X"13050d00",
		16#3ea0# => X"ef20103b",
		16#3ea1# => X"2322a100",
		16#3ea2# => X"93050d00",
		16#3ea3# => X"13050a00",
		16#3ea4# => X"ef20103a",
		16#3ea5# => X"2320a100",
		16#3ea6# => X"93850400",
		16#3ea7# => X"13050a00",
		16#3ea8# => X"ef201039",
		16#3ea9# => X"03284100",
		16#3eaa# => X"03278100",
		16#3eab# => X"83260100",
		16#3eac# => X"33050501",
		16#3ead# => X"93570701",
		16#3eae# => X"3385a700",
		16#3eaf# => X"63760501",
		16#3eb0# => X"0326c100",
		16#3eb1# => X"b386c600",
		16#3eb2# => X"93570501",
		16#3eb3# => X"37060100",
		16#3eb4# => X"b387d700",
		16#3eb5# => X"2320f102",
		16#3eb6# => X"9307f6ff",
		16#3eb7# => X"3375f500",
		16#3eb8# => X"13150501",
		16#3eb9# => X"3377f700",
		16#3eba# => X"3307e500",
		16#3ebb# => X"2328e102",
		16#3ebc# => X"03278106",
		16#3ebd# => X"93850900",
		16#3ebe# => X"232ec102",
		16#3ebf# => X"b377f700",
		16#3ec0# => X"93560701",
		16#3ec1# => X"13850700",
		16#3ec2# => X"2320d100",
		16#3ec3# => X"2324f100",
		16#3ec4# => X"ef201032",
		16#3ec5# => X"83258100",
		16#3ec6# => X"232ca102",
		16#3ec7# => X"13850a00",
		16#3ec8# => X"ef201031",
		16#3ec9# => X"83250100",
		16#3eca# => X"2326a100",
		16#3ecb# => X"13850a00",
		16#3ecc# => X"ef201030",
		16#3ecd# => X"2322a100",
		16#3ece# => X"03250100",
		16#3ecf# => X"93850900",
		16#3ed0# => X"ef20102f",
		16#3ed1# => X"0328c100",
		16#3ed2# => X"03278103",
		16#3ed3# => X"83264100",
		16#3ed4# => X"33050501",
		16#3ed5# => X"93570701",
		16#3ed6# => X"3385a700",
		16#3ed7# => X"63760501",
		16#3ed8# => X"0326c103",
		16#3ed9# => X"b386c600",
		16#3eda# => X"37080100",
		16#3edb# => X"93570501",
		16#3edc# => X"b386d700",
		16#3edd# => X"9307f8ff",
		16#3ede# => X"3376f500",
		16#3edf# => X"3377f700",
		16#3ee0# => X"13160601",
		16#3ee1# => X"3306e600",
		16#3ee2# => X"03278105",
		16#3ee3# => X"2326d104",
		16#3ee4# => X"93050400",
		16#3ee5# => X"b377f700",
		16#3ee6# => X"93560701",
		16#3ee7# => X"13850700",
		16#3ee8# => X"2322c104",
		16#3ee9# => X"2322d100",
		16#3eea# => X"2326f100",
		16#3eeb# => X"23240105",
		16#3eec# => X"ef201028",
		16#3eed# => X"2320a104",
		16#3eee# => X"03254100",
		16#3eef# => X"93050400",
		16#3ef0# => X"ef201027",
		16#3ef1# => X"83254100",
		16#3ef2# => X"232ea102",
		16#3ef3# => X"13050900",
		16#3ef4# => X"ef201026",
		16#3ef5# => X"8325c100",
		16#3ef6# => X"232ca102",
		16#3ef7# => X"13050900",
		16#3ef8# => X"ef201025",
		16#3ef9# => X"8328c103",
		16#3efa# => X"03230104",
		16#3efb# => X"03278103",
		16#3efc# => X"33051501",
		16#3efd# => X"93570301",
		16#3efe# => X"b387a700",
		16#3eff# => X"03264104",
		16#3f00# => X"8326c104",
		16#3f01# => X"63f61701",
		16#3f02# => X"03288104",
		16#3f03# => X"33070701",
		16#3f04# => X"13d80701",
		16#3f05# => X"3308e800",
		16#3f06# => X"37070100",
		16#3f07# => X"9305f7ff",
		16#3f08# => X"b3f7b700",
		16#3f09# => X"3373b300",
		16#3f0a# => X"93970701",
		16#3f0b# => X"b38e6700",
		16#3f0c# => X"83274103",
		16#3f0d# => X"232ce102",
		16#3f0e# => X"03270103",
		16#3f0f# => X"b38bfb00",
		16#3f10# => X"83278101",
		16#3f11# => X"b3bdbb01",
		16#3f12# => X"b388b701",
		16#3f13# => X"b3876b01",
		16#3f14# => X"33bb6701",
		16#3f15# => X"232cf100",
		16#3f16# => X"2322f108",
		16#3f17# => X"8327c101",
		16#3f18# => X"b3888801",
		16#3f19# => X"b387f800",
		16#3f1a# => X"338c6701",
		16#3f1b# => X"3303ec00",
		16#3f1c# => X"333ee300",
		16#3f1d# => X"0327c101",
		16#3f1e# => X"333c6c01",
		16#3f1f# => X"b3b8b801",
		16#3f20# => X"b3b7e700",
		16#3f21# => X"33ec8701",
		16#3f22# => X"83270102",
		16#3f23# => X"330c1c01",
		16#3f24# => X"3303c300",
		16#3f25# => X"330cfc00",
		16#3f26# => X"3305cc01",
		16#3f27# => X"b308d500",
		16#3f28# => X"03270102",
		16#3f29# => X"3336c300",
		16#3f2a# => X"b307d301",
		16#3f2b# => X"338fc800",
		16#3f2c# => X"33b3d701",
		16#3f2d# => X"232ef100",
		16#3f2e# => X"2324f108",
		16#3f2f# => X"032bc106",
		16#3f30# => X"b3070f01",
		16#3f31# => X"333ec501",
		16#3f32# => X"333cec00",
		16#3f33# => X"b3b6d800",
		16#3f34# => X"3336cf00",
		16#3f35# => X"b38d6700",
		16#3f36# => X"b3e6c600",
		16#3f37# => X"336ccc01",
		16#3f38# => X"b3b70701",
		16#3f39# => X"33b36d00",
		16#3f3a# => X"330cdc00",
		16#3f3b# => X"b3e76700",
		16#3f3c# => X"935b0b01",
		16#3f3d# => X"337bbb00",
		16#3f3e# => X"b307fc00",
		16#3f3f# => X"93850900",
		16#3f40# => X"13050b00",
		16#3f41# => X"2320f102",
		16#3f42# => X"ef209012",
		16#3f43# => X"130c0500",
		16#3f44# => X"93050b00",
		16#3f45# => X"13850a00",
		16#3f46# => X"ef209011",
		16#3f47# => X"2328a102",
		16#3f48# => X"93850b00",
		16#3f49# => X"13850a00",
		16#3f4a# => X"ef209010",
		16#3f4b# => X"930a0500",
		16#3f4c# => X"93850900",
		16#3f4d# => X"13850b00",
		16#3f4e# => X"ef20900f",
		16#3f4f# => X"83260103",
		16#3f50# => X"93570c01",
		16#3f51# => X"3305d500",
		16#3f52# => X"3385a700",
		16#3f53# => X"6376d500",
		16#3f54# => X"03278103",
		16#3f55# => X"b38aea00",
		16#3f56# => X"93570501",
		16#3f57# => X"b7060100",
		16#3f58# => X"b3875701",
		16#3f59# => X"2328f102",
		16#3f5a# => X"832ac105",
		16#3f5b# => X"9387f6ff",
		16#3f5c# => X"b379f500",
		16#3f5d# => X"337cfc00",
		16#3f5e# => X"93990901",
		16#3f5f# => X"b3898901",
		16#3f60# => X"13dc0a01",
		16#3f61# => X"b3fafa00",
		16#3f62# => X"93850a00",
		16#3f63# => X"13050400",
		16#3f64# => X"232ed102",
		16#3f65# => X"ef20d009",
		16#3f66# => X"93050400",
		16#3f67# => X"232ca102",
		16#3f68# => X"13050c00",
		16#3f69# => X"ef20d008",
		16#3f6a# => X"232aa102",
		16#3f6b# => X"93050c00",
		16#3f6c# => X"13050900",
		16#3f6d# => X"ef20d007",
		16#3f6e# => X"13040500",
		16#3f6f# => X"93850a00",
		16#3f70# => X"13050900",
		16#3f71# => X"ef20d006",
		16#3f72# => X"03264103",
		16#3f73# => X"03278103",
		16#3f74# => X"3305c500",
		16#3f75# => X"93570701",
		16#3f76# => X"3385a700",
		16#3f77# => X"6376c500",
		16#3f78# => X"8326c103",
		16#3f79# => X"3304d400",
		16#3f7a# => X"37080100",
		16#3f7b# => X"93570501",
		16#3f7c# => X"33848700",
		16#3f7d# => X"9307f8ff",
		16#3f7e# => X"3379f500",
		16#3f7f# => X"03258100",
		16#3f80# => X"3377f700",
		16#3f81# => X"93850400",
		16#3f82# => X"13190901",
		16#3f83# => X"23200105",
		16#3f84# => X"3309e900",
		16#3f85# => X"ef20d001",
		16#3f86# => X"83258100",
		16#3f87# => X"232ea102",
		16#3f88# => X"13050d00",
		16#3f89# => X"ef20d000",
		16#3f8a# => X"83250100",
		16#3f8b# => X"232ca102",
		16#3f8c# => X"13050d00",
		16#3f8d# => X"ef20c07f",
		16#3f8e# => X"232aa102",
		16#3f8f# => X"03250100",
		16#3f90# => X"93850400",
		16#3f91# => X"ef20c07e",
		16#3f92# => X"83288103",
		16#3f93# => X"8326c103",
		16#3f94# => X"03264103",
		16#3f95# => X"33051501",
		16#3f96# => X"93d70601",
		16#3f97# => X"3385a700",
		16#3f98# => X"63761501",
		16#3f99# => X"03280104",
		16#3f9a# => X"33060601",
		16#3f9b# => X"b7080100",
		16#3f9c# => X"9387f8ff",
		16#3f9d# => X"3377f500",
		16#3f9e# => X"135e0501",
		16#3f9f# => X"0325c100",
		16#3fa0# => X"b3f6f600",
		16#3fa1# => X"13170701",
		16#3fa2# => X"330ece00",
		16#3fa3# => X"3307d700",
		16#3fa4# => X"93850c00",
		16#3fa5# => X"2324c105",
		16#3fa6# => X"2320e104",
		16#3fa7# => X"23221105",
		16#3fa8# => X"ef200079",
		16#3fa9# => X"232ea102",
		16#3faa# => X"03254100",
		16#3fab# => X"93850c00",
		16#3fac# => X"ef200078",
		16#3fad# => X"83254100",
		16#3fae# => X"232ca102",
		16#3faf# => X"13050a00",
		16#3fb0# => X"ef200077",
		16#3fb1# => X"8325c100",
		16#3fb2# => X"232aa102",
		16#3fb3# => X"13050a00",
		16#3fb4# => X"ef200076",
		16#3fb5# => X"03238103",
		16#3fb6# => X"0328c103",
		16#3fb7# => X"03264103",
		16#3fb8# => X"33056500",
		16#3fb9# => X"93560801",
		16#3fba# => X"3385a600",
		16#3fbb# => X"03270104",
		16#3fbc# => X"032e8104",
		16#3fbd# => X"63766500",
		16#3fbe# => X"83284104",
		16#3fbf# => X"33061601",
		16#3fc0# => X"37030100",
		16#3fc1# => X"9306f3ff",
		16#3fc2# => X"93580501",
		16#3fc3# => X"b388c800",
		16#3fc4# => X"b377d500",
		16#3fc5# => X"3378d800",
		16#3fc6# => X"03260103",
		16#3fc7# => X"83260102",
		16#3fc8# => X"b38d3d01",
		16#3fc9# => X"b3bf3d01",
		16#3fca# => X"b386c600",
		16#3fcb# => X"338ff601",
		16#3fcc# => X"b38d2d01",
		16#3fcd# => X"93970701",
		16#3fce# => X"b3870701",
		16#3fcf# => X"33b92d01",
		16#3fd0# => X"33088f00",
		16#3fd1# => X"b30e2801",
		16#3fd2# => X"b38ded00",
		16#3fd3# => X"232a6102",
		16#3fd4# => X"03230103",
		16#3fd5# => X"b385ce01",
		16#3fd6# => X"33b7ed00",
		16#3fd7# => X"3386fd00",
		16#3fd8# => X"3385e500",
		16#3fd9# => X"33b92e01",
		16#3fda# => X"b3b5c501",
		16#3fdb# => X"b3b66600",
		16#3fdc# => X"333fff01",
		16#3fdd# => X"33348800",
		16#3fde# => X"b337f600",
		16#3fdf# => X"2320c102",
		16#3fe0# => X"2326c108",
		16#3fe1# => X"3337e500",
		16#3fe2# => X"33061501",
		16#3fe3# => X"33e7e500",
		16#3fe4# => X"33efe601",
		16#3fe5# => X"b309f600",
		16#3fe6# => X"33642401",
		16#3fe7# => X"8325c100",
		16#3fe8# => X"03258100",
		16#3fe9# => X"33048f00",
		16#3fea# => X"33361601",
		16#3feb# => X"b3b7f900",
		16#3fec# => X"3304e400",
		16#3fed# => X"b367f600",
		16#3fee# => X"3304f400",
		16#3fef# => X"ef204067",
		16#3ff0# => X"2328a102",
		16#3ff1# => X"83258100",
		16#3ff2# => X"03254100",
		16#3ff3# => X"ef204066",
		16#3ff4# => X"13090500",
		16#3ff5# => X"83254100",
		16#3ff6# => X"03250100",
		16#3ff7# => X"ef204065",
		16#3ff8# => X"930d0500",
		16#3ff9# => X"8325c100",
		16#3ffa# => X"03250100",
		16#3ffb# => X"ef204064",
		16#3ffc# => X"03270103",
		16#3ffd# => X"33052501",
		16#3ffe# => X"93570701",
		16#3fff# => X"3385a700",
		16#4000# => X"63762501",
		16#4001# => X"03234103",
		16#4002# => X"b38d6d00",
		16#4003# => X"b7060100",
		16#4004# => X"93570501",
		16#4005# => X"b38db701",
		16#4006# => X"9387f6ff",
		16#4007# => X"3379f500",
		16#4008# => X"3377f700",
		16#4009# => X"93850400",
		16#400a# => X"13190901",
		16#400b# => X"13050b00",
		16#400c# => X"3309e900",
		16#400d# => X"232cd102",
		16#400e# => X"ef20805f",
		16#400f# => X"232aa102",
		16#4010# => X"93050b00",
		16#4011# => X"13050d00",
		16#4012# => X"ef20805e",
		16#4013# => X"2328a102",
		16#4014# => X"93850b00",
		16#4015# => X"13050d00",
		16#4016# => X"ef20805d",
		16#4017# => X"130d0500",
		16#4018# => X"93850400",
		16#4019# => X"13850b00",
		16#401a# => X"ef20805c",
		16#401b# => X"03260103",
		16#401c# => X"03274103",
		16#401d# => X"3305c500",
		16#401e# => X"93570701",
		16#401f# => X"3385a700",
		16#4020# => X"6376c500",
		16#4021# => X"83268103",
		16#4022# => X"330ddd00",
		16#4023# => X"b7060100",
		16#4024# => X"93570501",
		16#4025# => X"338da701",
		16#4026# => X"9387f6ff",
		16#4027# => X"b374f500",
		16#4028# => X"3377f700",
		16#4029# => X"93850c00",
		16#402a# => X"93940401",
		16#402b# => X"13850a00",
		16#402c# => X"b384e400",
		16#402d# => X"232cd102",
		16#402e# => X"ef208057",
		16#402f# => X"93850c00",
		16#4030# => X"232aa102",
		16#4031# => X"13050c00",
		16#4032# => X"ef208056",
		16#4033# => X"2328a102",
		16#4034# => X"93050c00",
		16#4035# => X"13050a00",
		16#4036# => X"ef208055",
		16#4037# => X"930c0500",
		16#4038# => X"93850a00",
		16#4039# => X"13050a00",
		16#403a# => X"ef208054",
		16#403b# => X"03260103",
		16#403c# => X"03274103",
		16#403d# => X"3305c500",
		16#403e# => X"93570701",
		16#403f# => X"3385a700",
		16#4040# => X"6376c500",
		16#4041# => X"83268103",
		16#4042# => X"b38cdc00",
		16#4043# => X"37080100",
		16#4044# => X"93570501",
		16#4045# => X"b38c9701",
		16#4046# => X"9307f8ff",
		16#4047# => X"337af500",
		16#4048# => X"0325c100",
		16#4049# => X"3377f700",
		16#404a# => X"93050b00",
		16#404b# => X"131a0a01",
		16#404c# => X"330aea00",
		16#404d# => X"232c0103",
		16#404e# => X"ef20804f",
		16#404f# => X"232aa102",
		16#4050# => X"03254100",
		16#4051# => X"93050b00",
		16#4052# => X"ef20804e",
		16#4053# => X"2328a102",
		16#4054# => X"03254100",
		16#4055# => X"93850b00",
		16#4056# => X"ef20804d",
		16#4057# => X"8325c100",
		16#4058# => X"2322a100",
		16#4059# => X"13850b00",
		16#405a# => X"ef20804c",
		16#405b# => X"83280103",
		16#405c# => X"83264103",
		16#405d# => X"03264100",
		16#405e# => X"33051501",
		16#405f# => X"13d70601",
		16#4060# => X"3305a700",
		16#4061# => X"63761501",
		16#4062# => X"03288103",
		16#4063# => X"33060601",
		16#4064# => X"37080100",
		16#4065# => X"1307f8ff",
		16#4066# => X"b377e500",
		16#4067# => X"13530501",
		16#4068# => X"03258100",
		16#4069# => X"b3f6e600",
		16#406a# => X"93970701",
		16#406b# => X"3303c300",
		16#406c# => X"b387d700",
		16#406d# => X"93850a00",
		16#406e# => X"232c6102",
		16#406f# => X"2328f102",
		16#4070# => X"232a0103",
		16#4071# => X"ef20c046",
		16#4072# => X"83258100",
		16#4073# => X"2326a100",
		16#4074# => X"13050c00",
		16#4075# => X"ef20c045",
		16#4076# => X"2324a100",
		16#4077# => X"03250100",
		16#4078# => X"93050c00",
		16#4079# => X"ef20c044",
		16#407a# => X"2322a100",
		16#407b# => X"03250100",
		16#407c# => X"93850a00",
		16#407d# => X"ef20c043",
		16#407e# => X"83288100",
		16#407f# => X"032ec100",
		16#4080# => X"03264100",
		16#4081# => X"33051501",
		16#4082# => X"93560e01",
		16#4083# => X"3385a600",
		16#4084# => X"83270103",
		16#4085# => X"03238103",
		16#4086# => X"63761501",
		16#4087# => X"03284103",
		16#4088# => X"33060601",
		16#4089# => X"37080100",
		16#408a# => X"93580501",
		16#408b# => X"b3892901",
		16#408c# => X"b388c800",
		16#408d# => X"33b92901",
		16#408e# => X"1306f8ff",
		16#408f# => X"3304b401",
		16#4090# => X"b30e2401",
		16#4091# => X"3377c500",
		16#4092# => X"b3899900",
		16#4093# => X"337ece00",
		16#4094# => X"b385ae01",
		16#4095# => X"b3b49900",
		16#4096# => X"13170701",
		16#4097# => X"3307c701",
		16#4098# => X"b3894901",
		16#4099# => X"338e9500",
		16#409a# => X"330f9e01",
		16#409b# => X"33ba4901",
		16#409c# => X"b30f4f01",
		16#409d# => X"33b52e01",
		16#409e# => X"3334b401",
		16#409f# => X"33bda501",
		16#40a0# => X"b3349e00",
		16#40a1# => X"336e9d00",
		16#40a2# => X"b33c9f01",
		16#40a3# => X"33ba4f01",
		16#40a4# => X"3365a400",
		16#40a5# => X"3305c501",
		16#40a6# => X"33ea4c01",
		16#40a7# => X"b386ff00",
		16#40a8# => X"33054501",
		16#40a9# => X"33056500",
		16#40aa# => X"b3b7f600",
		16#40ab# => X"b305f500",
		16#40ac# => X"b3b7f500",
		16#40ad# => X"33356500",
		16#40ae# => X"b386e600",
		16#40af# => X"33b7e600",
		16#40b0# => X"3364f500",
		16#40b1# => X"33851501",
		16#40b2# => X"b304e500",
		16#40b3# => X"33b7e400",
		16#40b4# => X"33351501",
		16#40b5# => X"23283109",
		16#40b6# => X"93850a00",
		16#40b7# => X"b369e500",
		16#40b8# => X"13050b00",
		16#40b9# => X"2320c100",
		16#40ba# => X"23220101",
		16#40bb# => X"232ad108",
		16#40bc# => X"ef200034",
		16#40bd# => X"93050b00",
		16#40be# => X"130a0500",
		16#40bf# => X"13050c00",
		16#40c0# => X"ef200033",
		16#40c1# => X"130b0500",
		16#40c2# => X"93050c00",
		16#40c3# => X"13850b00",
		16#40c4# => X"ef200032",
		16#40c5# => X"13090500",
		16#40c6# => X"93850a00",
		16#40c7# => X"13850b00",
		16#40c8# => X"ef200031",
		16#40c9# => X"33056501",
		16#40ca# => X"13570a01",
		16#40cb# => X"3305a700",
		16#40cc# => X"03260100",
		16#40cd# => X"63766501",
		16#40ce# => X"03284100",
		16#40cf# => X"33090901",
		16#40d0# => X"b377c500",
		16#40d1# => X"93970701",
		16#40d2# => X"3376ca00",
		16#40d3# => X"3386c700",
		16#40d4# => X"03278101",
		16#40d5# => X"8327c102",
		16#40d6# => X"13550501",
		16#40d7# => X"b384c400",
		16#40d8# => X"b3e7e700",
		16#40d9# => X"0327c101",
		16#40da# => X"33058500",
		16#40db# => X"33b6c400",
		16#40dc# => X"b36bf700",
		16#40dd# => X"83270102",
		16#40de# => X"33053501",
		16#40df# => X"3305c500",
		16#40e0# => X"33052501",
		16#40e1# => X"9397d700",
		16#40e2# => X"232ea108",
		16#40e3# => X"232c9108",
		16#40e4# => X"b3e77701",
		16#40e5# => X"13070108",
		16#40e6# => X"13060000",
		16#40e7# => X"13054000",
		16#40e8# => X"8326c700",
		16#40e9# => X"83250701",
		16#40ea# => X"13061600",
		16#40eb# => X"93d63601",
		16#40ec# => X"9395d500",
		16#40ed# => X"b3e6b600",
		16#40ee# => X"2320d700",
		16#40ef# => X"13074700",
		16#40f0# => X"e310a6fe",
		16#40f1# => X"03270108",
		16#40f2# => X"83268108",
		16#40f3# => X"b337f000",
		16#40f4# => X"b3e7e700",
		16#40f5# => X"232cd106",
		16#40f6# => X"0327c108",
		16#40f7# => X"83264108",
		16#40f8# => X"2328f106",
		16#40f9# => X"232ee106",
		16#40fa# => X"232ad106",
		16#40fb# => X"9316b700",
		16#40fc# => X"63d40624",
		16#40fd# => X"9397f701",
		16#40fe# => X"13070107",
		16#40ff# => X"13060000",
		16#4100# => X"13053000",
		16#4101# => X"83260700",
		16#4102# => X"83254700",
		16#4103# => X"13061600",
		16#4104# => X"93d61600",
		16#4105# => X"9395f501",
		16#4106# => X"b3e6b600",
		16#4107# => X"2320d700",
		16#4108# => X"13074700",
		16#4109# => X"e310a6fe",
		16#410a# => X"0327c107",
		16#410b# => X"b337f000",
		16#410c# => X"13571700",
		16#410d# => X"232ee106",
		16#410e# => X"03270107",
		16#410f# => X"b367f700",
		16#4110# => X"2328f106",
		16#4111# => X"03274102",
		16#4112# => X"b7470000",
		16#4113# => X"9387f7ff",
		16#4114# => X"b307f700",
		16#4115# => X"6354f020",
		16#4116# => X"03270107",
		16#4117# => X"93767700",
		16#4118# => X"63840604",
		16#4119# => X"9376f700",
		16#411a# => X"13064000",
		16#411b# => X"638ec602",
		16#411c# => X"83264107",
		16#411d# => X"13074700",
		16#411e# => X"2328e106",
		16#411f# => X"13374700",
		16#4120# => X"b306d700",
		16#4121# => X"33b7e600",
		16#4122# => X"232ad106",
		16#4123# => X"83268107",
		16#4124# => X"b306d700",
		16#4125# => X"232cd106",
		16#4126# => X"b3b6e600",
		16#4127# => X"0327c107",
		16#4128# => X"b386e600",
		16#4129# => X"232ed106",
		16#412a# => X"0327c107",
		16#412b# => X"9316b700",
		16#412c# => X"63d00602",
		16#412d# => X"b707f0ff",
		16#412e# => X"9387f7ff",
		16#412f# => X"3377f700",
		16#4130# => X"232ee106",
		16#4131# => X"03274102",
		16#4132# => X"b7470000",
		16#4133# => X"b307f700",
		16#4134# => X"13070107",
		16#4135# => X"13060000",
		16#4136# => X"13053000",
		16#4137# => X"83260700",
		16#4138# => X"83254700",
		16#4139# => X"13061600",
		16#413a# => X"93d63600",
		16#413b# => X"9395d501",
		16#413c# => X"b3e6b600",
		16#413d# => X"2320d700",
		16#413e# => X"13074700",
		16#413f# => X"e310a6fe",
		16#4140# => X"37870000",
		16#4141# => X"9306e7ff",
		16#4142# => X"63cef612",
		16#4143# => X"0327c107",
		16#4144# => X"13573700",
		16#4145# => X"232ee106",
		16#4146# => X"0327c107",
		16#4147# => X"b7060180",
		16#4148# => X"9386f6ff",
		16#4149# => X"2316e108",
		16#414a# => X"37870000",
		16#414b# => X"1307f7ff",
		16#414c# => X"b3f7e700",
		16#414d# => X"0327c108",
		16#414e# => X"93970701",
		16#414f# => X"8320c10d",
		16#4150# => X"3377d700",
		16#4151# => X"b367f700",
		16#4152# => X"03274101",
		16#4153# => X"b7060080",
		16#4154# => X"93c6f6ff",
		16#4155# => X"1317f701",
		16#4156# => X"b3f7d700",
		16#4157# => X"b3e7e700",
		16#4158# => X"83260101",
		16#4159# => X"03270107",
		16#415a# => X"0324810d",
		16#415b# => X"23a6f600",
		16#415c# => X"23a0e600",
		16#415d# => X"03274107",
		16#415e# => X"8324410d",
		16#415f# => X"0329010d",
		16#4160# => X"23a2e600",
		16#4161# => X"03278107",
		16#4162# => X"8329c10c",
		16#4163# => X"032a810c",
		16#4164# => X"23a4e600",
		16#4165# => X"832a410c",
		16#4166# => X"032b010c",
		16#4167# => X"832bc10b",
		16#4168# => X"032c810b",
		16#4169# => X"832c410b",
		16#416a# => X"032d010b",
		16#416b# => X"832dc10a",
		16#416c# => X"13850600",
		16#416d# => X"1301010e",
		16#416e# => X"67800000",
		16#416f# => X"232a3101",
		16#4170# => X"83270105",
		16#4171# => X"2328f106",
		16#4172# => X"83274105",
		16#4173# => X"232af106",
		16#4174# => X"83278105",
		16#4175# => X"232cf106",
		16#4176# => X"8327c105",
		16#4177# => X"232ef106",
		16#4178# => X"93072000",
		16#4179# => X"6380f428",
		16#417a# => X"93073000",
		16#417b# => X"638af428",
		16#417c# => X"93071000",
		16#417d# => X"e398f4e4",
		16#417e# => X"232e0106",
		16#417f# => X"232c0106",
		16#4180# => X"232a0106",
		16#4181# => X"23280106",
		16#4182# => X"6f00c021",
		16#4183# => X"232a2101",
		16#4184# => X"83270106",
		16#4185# => X"93040700",
		16#4186# => X"2328f106",
		16#4187# => X"83274106",
		16#4188# => X"232af106",
		16#4189# => X"83278106",
		16#418a# => X"232cf106",
		16#418b# => X"8327c106",
		16#418c# => X"232ef106",
		16#418d# => X"6ff0dffa",
		16#418e# => X"83278102",
		16#418f# => X"2322f102",
		16#4190# => X"6ff05fe0",
		16#4191# => X"232e0106",
		16#4192# => X"232c0106",
		16#4193# => X"232a0106",
		16#4194# => X"23280106",
		16#4195# => X"9307f7ff",
		16#4196# => X"6ff01fec",
		16#4197# => X"93061000",
		16#4198# => X"b387f640",
		16#4199# => X"13074007",
		16#419a# => X"6342f71c",
		16#419b# => X"13d65740",
		16#419c# => X"93f6f701",
		16#419d# => X"13070000",
		16#419e# => X"93070000",
		16#419f# => X"93152700",
		16#41a0# => X"6312c702",
		16#41a1# => X"63980604",
		16#41a2# => X"13053000",
		16#41a3# => X"13060107",
		16#41a4# => X"3305e540",
		16#41a5# => X"6354d502",
		16#41a6# => X"93064000",
		16#41a7# => X"3387e640",
		16#41a8# => X"6f004008",
		16#41a9# => X"13050107",
		16#41aa# => X"b305b500",
		16#41ab# => X"83a50500",
		16#41ac# => X"13071700",
		16#41ad# => X"b3e7b700",
		16#41ae# => X"6ff05ffc",
		16#41af# => X"3308b600",
		16#41b0# => X"03280800",
		16#41b1# => X"93861600",
		16#41b2# => X"13064600",
		16#41b3# => X"232e06ff",
		16#41b4# => X"6ff05ffc",
		16#41b5# => X"1306010a",
		16#41b6# => X"3306b600",
		16#41b7# => X"032606fd",
		16#41b8# => X"13080002",
		16#41b9# => X"3308d840",
		16#41ba# => X"33160601",
		16#41bb# => X"b3e7c700",
		16#41bc# => X"13063000",
		16#41bd# => X"93080107",
		16#41be# => X"13030000",
		16#41bf# => X"3306e640",
		16#41c0# => X"6346c302",
		16#41c1# => X"93054000",
		16#41c2# => X"3387e540",
		16#41c3# => X"13162600",
		16#41c4# => X"9305010a",
		16#41c5# => X"3386c500",
		16#41c6# => X"8325c107",
		16#41c7# => X"b3d6d500",
		16#41c8# => X"2328d6fc",
		16#41c9# => X"13064000",
		16#41ca# => X"6f000004",
		16#41cb# => X"338eb800",
		16#41cc# => X"03250e00",
		16#41cd# => X"032e4e00",
		16#41ce# => X"13031300",
		16#41cf# => X"3355d500",
		16#41d0# => X"331e0e01",
		16#41d1# => X"3365c501",
		16#41d2# => X"23a0a800",
		16#41d3# => X"93884800",
		16#41d4# => X"6ff01ffb",
		16#41d5# => X"93162700",
		16#41d6# => X"93050107",
		16#41d7# => X"b386d500",
		16#41d8# => X"23a00600",
		16#41d9# => X"13071700",
		16#41da# => X"e316c7fe",
		16#41db# => X"83260107",
		16#41dc# => X"b337f000",
		16#41dd# => X"b3e7d700",
		16#41de# => X"2328f106",
		16#41df# => X"93f67700",
		16#41e0# => X"63820604",
		16#41e1# => X"93f6f700",
		16#41e2# => X"638ee602",
		16#41e3# => X"03274107",
		16#41e4# => X"93874700",
		16#41e5# => X"2328f106",
		16#41e6# => X"93b74700",
		16#41e7# => X"3387e700",
		16#41e8# => X"b337f700",
		16#41e9# => X"232ae106",
		16#41ea# => X"03278107",
		16#41eb# => X"3387e700",
		16#41ec# => X"232ce106",
		16#41ed# => X"3337f700",
		16#41ee# => X"8327c107",
		16#41ef# => X"3307f700",
		16#41f0# => X"232ee106",
		16#41f1# => X"8327c107",
		16#41f2# => X"1397c700",
		16#41f3# => X"635e0700",
		16#41f4# => X"232e0106",
		16#41f5# => X"232c0106",
		16#41f6# => X"232a0106",
		16#41f7# => X"23280106",
		16#41f8# => X"93071000",
		16#41f9# => X"6ff05fd3",
		16#41fa# => X"93070107",
		16#41fb# => X"93060000",
		16#41fc# => X"93053000",
		16#41fd# => X"03a70700",
		16#41fe# => X"03a64700",
		16#41ff# => X"93861600",
		16#4200# => X"13573700",
		16#4201# => X"1316d601",
		16#4202# => X"3367c700",
		16#4203# => X"23a0e700",
		16#4204# => X"93874700",
		16#4205# => X"e390b6fe",
		16#4206# => X"8327c107",
		16#4207# => X"93d73700",
		16#4208# => X"232ef106",
		16#4209# => X"93070000",
		16#420a# => X"6ff01fcf",
		16#420b# => X"83274107",
		16#420c# => X"03270107",
		16#420d# => X"3367f700",
		16#420e# => X"83278107",
		16#420f# => X"3367f700",
		16#4210# => X"8327c107",
		16#4211# => X"3367f700",
		16#4212# => X"93070000",
		16#4213# => X"e30607cc",
		16#4214# => X"232e0106",
		16#4215# => X"232c0106",
		16#4216# => X"232a0106",
		16#4217# => X"23280106",
		16#4218# => X"6ff09fcb",
		16#4219# => X"b7870000",
		16#421a# => X"232e0106",
		16#421b# => X"232c0106",
		16#421c# => X"232a0106",
		16#421d# => X"23280106",
		16#421e# => X"9387f7ff",
		16#421f# => X"6ff0dfc9",
		16#4220# => X"b7870000",
		16#4221# => X"232ef106",
		16#4222# => X"232c0106",
		16#4223# => X"232a0106",
		16#4224# => X"23280106",
		16#4225# => X"9387f7ff",
		16#4226# => X"232a0100",
		16#4227# => X"6ff0dfc7",
		16#4228# => X"130101fa",
		16#4229# => X"83a78500",
		16#422a# => X"23244105",
		16#422b# => X"03aac500",
		16#422c# => X"83a60500",
		16#422d# => X"03a74500",
		16#422e# => X"232cf102",
		16#422f# => X"232cf100",
		16#4230# => X"93170a01",
		16#4231# => X"232c8104",
		16#4232# => X"93d70701",
		16#4233# => X"13141a00",
		16#4234# => X"232a9104",
		16#4235# => X"03230600",
		16#4236# => X"93040500",
		16#4237# => X"83284600",
		16#4238# => X"83258600",
		16#4239# => X"0325c600",
		16#423a# => X"232e4103",
		16#423b# => X"232e1104",
		16#423c# => X"23282105",
		16#423d# => X"23263105",
		16#423e# => X"23225105",
		16#423f# => X"2328d102",
		16#4240# => X"232ae102",
		16#4241# => X"2328d100",
		16#4242# => X"232ae100",
		16#4243# => X"232ef100",
		16#4244# => X"13541401",
		16#4245# => X"135afa01",
		16#4246# => X"13080101",
		16#4247# => X"1306c101",
		16#4248# => X"83270600",
		16#4249# => X"0327c6ff",
		16#424a# => X"1306c6ff",
		16#424b# => X"93973700",
		16#424c# => X"1357d701",
		16#424d# => X"b3e7e700",
		16#424e# => X"2322f600",
		16#424f# => X"e312c8fe",
		16#4250# => X"83260101",
		16#4251# => X"93170501",
		16#4252# => X"232cb102",
		16#4253# => X"93963600",
		16#4254# => X"2324b102",
		16#4255# => X"93d70701",
		16#4256# => X"93151500",
		16#4257# => X"23286102",
		16#4258# => X"232a1103",
		16#4259# => X"232ea102",
		16#425a# => X"23206102",
		16#425b# => X"23221103",
		16#425c# => X"2328d100",
		16#425d# => X"2326f102",
		16#425e# => X"93d51501",
		16#425f# => X"1355f501",
		16#4260# => X"93080102",
		16#4261# => X"1303c102",
		16#4262# => X"83270300",
		16#4263# => X"0327c3ff",
		16#4264# => X"1303c3ff",
		16#4265# => X"93973700",
		16#4266# => X"1357d701",
		16#4267# => X"b3e7e700",
		16#4268# => X"2322f300",
		16#4269# => X"e39268fe",
		16#426a# => X"83270102",
		16#426b# => X"37870000",
		16#426c# => X"1307f7ff",
		16#426d# => X"93973700",
		16#426e# => X"2320f102",
		16#426f# => X"6390e502",
		16#4270# => X"032e8102",
		16#4271# => X"03274102",
		16#4272# => X"3367c701",
		16#4273# => X"032ec102",
		16#4274# => X"3367c701",
		16#4275# => X"3367f700",
		16#4276# => X"63140700",
		16#4277# => X"13451500",
		16#4278# => X"3307b440",
		16#4279# => X"e3164511",
		16#427a# => X"6352e030",
		16#427b# => X"63960514",
		16#427c# => X"03254102",
		16#427d# => X"83258102",
		16#427e# => X"0328c102",
		16#427f# => X"3366b500",
		16#4280# => X"33660601",
		16#4281# => X"3366f600",
		16#4282# => X"63140602",
		16#4283# => X"83274101",
		16#4284# => X"2328d102",
		16#4285# => X"13040700",
		16#4286# => X"232af102",
		16#4287# => X"83278101",
		16#4288# => X"232cf102",
		16#4289# => X"8327c101",
		16#428a# => X"232ef102",
		16#428b# => X"6f004030",
		16#428c# => X"1306f7ff",
		16#428d# => X"631e060c",
		16#428e# => X"03274101",
		16#428f# => X"b387f600",
		16#4290# => X"b3b6d700",
		16#4291# => X"3306e500",
		16#4292# => X"2328f102",
		16#4293# => X"b307d600",
		16#4294# => X"b3b6d700",
		16#4295# => X"232af102",
		16#4296# => X"83278101",
		16#4297# => X"3337e600",
		16#4298# => X"b366d700",
		16#4299# => X"3387f500",
		16#429a# => X"3306d700",
		16#429b# => X"b337f700",
		16#429c# => X"0327c101",
		16#429d# => X"b336d600",
		16#429e# => X"b3e7d700",
		16#429f# => X"3308e800",
		16#42a0# => X"b3870701",
		16#42a1# => X"232cc102",
		16#42a2# => X"232ef102",
		16#42a3# => X"13041000",
		16#42a4# => X"8327c103",
		16#42a5# => X"1397c700",
		16#42a6# => X"635c0728",
		16#42a7# => X"3707f8ff",
		16#42a8# => X"1307f7ff",
		16#42a9# => X"b3f7e700",
		16#42aa# => X"232ef102",
		16#42ab# => X"83270103",
		16#42ac# => X"13041400",
		16#42ad# => X"13070103",
		16#42ae# => X"9397f701",
		16#42af# => X"13060000",
		16#42b0# => X"13053000",
		16#42b1# => X"83260700",
		16#42b2# => X"83254700",
		16#42b3# => X"13061600",
		16#42b4# => X"93d61600",
		16#42b5# => X"9395f501",
		16#42b6# => X"b3e6b600",
		16#42b7# => X"2320d700",
		16#42b8# => X"13074700",
		16#42b9# => X"e310a6fe",
		16#42ba# => X"0327c103",
		16#42bb# => X"b337f000",
		16#42bc# => X"13571700",
		16#42bd# => X"232ee102",
		16#42be# => X"03270103",
		16#42bf# => X"b367f700",
		16#42c0# => X"2328f102",
		16#42c1# => X"b7870000",
		16#42c2# => X"9387f7ff",
		16#42c3# => X"6f00c07c",
		16#42c4# => X"b7870000",
		16#42c5# => X"9387f7ff",
		16#42c6# => X"e30af7ee",
		16#42c7# => X"93074007",
		16#42c8# => X"63d0c706",
		16#42c9# => X"23260102",
		16#42ca# => X"23240102",
		16#42cb# => X"23220102",
		16#42cc# => X"93071000",
		16#42cd# => X"6f008014",
		16#42ce# => X"b7870000",
		16#42cf# => X"9387f7ff",
		16#42d0# => X"6312f402",
		16#42d1# => X"83274101",
		16#42d2# => X"2328d102",
		16#42d3# => X"232af102",
		16#42d4# => X"83278101",
		16#42d5# => X"232cf102",
		16#42d6# => X"8327c101",
		16#42d7# => X"232ef102",
		16#42d8# => X"6f00001d",
		16#42d9# => X"8327c102",
		16#42da# => X"b7060800",
		16#42db# => X"b3e7d700",
		16#42dc# => X"2326f102",
		16#42dd# => X"93074007",
		16#42de# => X"e3c6e7fa",
		16#42df# => X"13060700",
		16#42e0# => X"13575640",
		16#42e1# => X"93050000",
		16#42e2# => X"1376f601",
		16#42e3# => X"93070000",
		16#42e4# => X"93962700",
		16#42e5# => X"6390e702",
		16#42e6# => X"63140604",
		16#42e7# => X"13073000",
		16#42e8# => X"3307f740",
		16#42e9# => X"6352c702",
		16#42ea# => X"13074000",
		16#42eb# => X"b307f740",
		16#42ec# => X"6f00c007",
		16#42ed# => X"b386d800",
		16#42ee# => X"83a60600",
		16#42ef# => X"93871700",
		16#42f0# => X"b3e5d500",
		16#42f1# => X"6ff0dffc",
		16#42f2# => X"3305d300",
		16#42f3# => X"03250500",
		16#42f4# => X"13061600",
		16#42f5# => X"13034300",
		16#42f6# => X"232ea3fe",
		16#42f7# => X"6ff09ffc",
		16#42f8# => X"13070104",
		16#42f9# => X"3307d700",
		16#42fa# => X"032707fe",
		16#42fb# => X"13080002",
		16#42fc# => X"3308c840",
		16#42fd# => X"33170701",
		16#42fe# => X"b3e5e500",
		16#42ff# => X"13073000",
		16#4300# => X"130e0000",
		16#4301# => X"3307f740",
		16#4302# => X"6346ee02",
		16#4303# => X"93064000",
		16#4304# => X"b387f640",
		16#4305# => X"13172700",
		16#4306# => X"93060104",
		16#4307# => X"3387e600",
		16#4308# => X"8326c102",
		16#4309# => X"33d6c600",
		16#430a# => X"2320c7fe",
		16#430b# => X"93064000",
		16#430c# => X"6f00c003",
		16#430d# => X"b30ed300",
		16#430e# => X"03a50e00",
		16#430f# => X"83ae4e00",
		16#4310# => X"130e1e00",
		16#4311# => X"3355c500",
		16#4312# => X"b39e0e01",
		16#4313# => X"3365d501",
		16#4314# => X"2320a300",
		16#4315# => X"13034300",
		16#4316# => X"6ff01ffb",
		16#4317# => X"13972700",
		16#4318# => X"3387e800",
		16#4319# => X"23200700",
		16#431a# => X"93871700",
		16#431b# => X"e398d7fe",
		16#431c# => X"03270102",
		16#431d# => X"b337b000",
		16#431e# => X"b367f700",
		16#431f# => X"2320f102",
		16#4320# => X"83260101",
		16#4321# => X"83270102",
		16#4322# => X"03274101",
		16#4323# => X"83258102",
		16#4324# => X"b387f600",
		16#4325# => X"b3b6d700",
		16#4326# => X"2328f102",
		16#4327# => X"83274102",
		16#4328# => X"0325c102",
		16#4329# => X"b307f700",
		16#432a# => X"3386d700",
		16#432b# => X"33b7e700",
		16#432c# => X"b337d600",
		16#432d# => X"b367f700",
		16#432e# => X"03278101",
		16#432f# => X"8326c101",
		16#4330# => X"232ac102",
		16#4331# => X"b305b700",
		16#4332# => X"3386f500",
		16#4333# => X"33b7e500",
		16#4334# => X"b337f600",
		16#4335# => X"b386a600",
		16#4336# => X"3367f700",
		16#4337# => X"3387e600",
		16#4338# => X"232cc102",
		16#4339# => X"232ee102",
		16#433a# => X"6ff09fda",
		16#433b# => X"6300073e",
		16#433c# => X"63160424",
		16#433d# => X"83284101",
		16#433e# => X"03258101",
		16#433f# => X"032ec101",
		16#4340# => X"33e3a800",
		16#4341# => X"3363c301",
		16#4342# => X"3363d300",
		16#4343# => X"6310031a",
		16#4344# => X"2328f102",
		16#4345# => X"83274102",
		16#4346# => X"13840500",
		16#4347# => X"232af102",
		16#4348# => X"83278102",
		16#4349# => X"232cf102",
		16#434a# => X"8327c102",
		16#434b# => X"232ef102",
		16#434c# => X"83270103",
		16#434d# => X"13f77700",
		16#434e# => X"63040704",
		16#434f# => X"13f7f700",
		16#4350# => X"93064000",
		16#4351# => X"630ed702",
		16#4352# => X"03274103",
		16#4353# => X"93874700",
		16#4354# => X"2328f102",
		16#4355# => X"93b74700",
		16#4356# => X"3387e700",
		16#4357# => X"b337f700",
		16#4358# => X"232ae102",
		16#4359# => X"03278103",
		16#435a# => X"3387e700",
		16#435b# => X"232ce102",
		16#435c# => X"3337f700",
		16#435d# => X"8327c103",
		16#435e# => X"3307f700",
		16#435f# => X"232ee102",
		16#4360# => X"8327c103",
		16#4361# => X"1397c700",
		16#4362# => X"63540702",
		16#4363# => X"37870000",
		16#4364# => X"13041400",
		16#4365# => X"1307f7ff",
		16#4366# => X"6314e400",
		16#4367# => X"6f00507f",
		16#4368# => X"3707f8ff",
		16#4369# => X"1307f7ff",
		16#436a# => X"b3f7e700",
		16#436b# => X"232ef102",
		16#436c# => X"93070103",
		16#436d# => X"93060000",
		16#436e# => X"93053000",
		16#436f# => X"03a70700",
		16#4370# => X"03a64700",
		16#4371# => X"93861600",
		16#4372# => X"13573700",
		16#4373# => X"1316d601",
		16#4374# => X"3367c700",
		16#4375# => X"23a0e700",
		16#4376# => X"93874700",
		16#4377# => X"e390b6fe",
		16#4378# => X"8327c103",
		16#4379# => X"b7860000",
		16#437a# => X"13d73700",
		16#437b# => X"232ee102",
		16#437c# => X"9387f6ff",
		16#437d# => X"631af402",
		16#437e# => X"03264103",
		16#437f# => X"83270103",
		16#4380# => X"b3e7c700",
		16#4381# => X"03268103",
		16#4382# => X"b3e7c700",
		16#4383# => X"b3e7e700",
		16#4384# => X"638c0700",
		16#4385# => X"232ed102",
		16#4386# => X"232c0102",
		16#4387# => X"232a0102",
		16#4388# => X"23280102",
		16#4389# => X"130a0000",
		16#438a# => X"8327c103",
		16#438b# => X"37070180",
		16#438c# => X"1307f7ff",
		16#438d# => X"2316f100",
		16#438e# => X"b7870000",
		16#438f# => X"9387f7ff",
		16#4390# => X"3374f400",
		16#4391# => X"93170401",
		16#4392# => X"0324c100",
		16#4393# => X"8320c105",
		16#4394# => X"13850400",
		16#4395# => X"3374e400",
		16#4396# => X"3364f400",
		16#4397# => X"9317fa01",
		16#4398# => X"370a0080",
		16#4399# => X"134afaff",
		16#439a# => X"33744401",
		16#439b# => X"336af400",
		16#439c# => X"83270103",
		16#439d# => X"03248105",
		16#439e# => X"23a64401",
		16#439f# => X"23a0f400",
		16#43a0# => X"83274103",
		16#43a1# => X"03290105",
		16#43a2# => X"8329c104",
		16#43a3# => X"23a2f400",
		16#43a4# => X"83278103",
		16#43a5# => X"032a8104",
		16#43a6# => X"832a4104",
		16#43a7# => X"23a4f400",
		16#43a8# => X"83244105",
		16#43a9# => X"13010106",
		16#43aa# => X"67800000",
		16#43ab# => X"1303f0ff",
		16#43ac# => X"63106706",
		16#43ad# => X"03264102",
		16#43ae# => X"b386f600",
		16#43af# => X"b3b7f600",
		16#43b0# => X"3388c800",
		16#43b1# => X"3307f800",
		16#43b2# => X"b337f700",
		16#43b3# => X"232ae102",
		16#43b4# => X"03278102",
		16#43b5# => X"3336c800",
		16#43b6# => X"b367f600",
		16#43b7# => X"2328d102",
		16#43b8# => X"b306e500",
		16#43b9# => X"3386f600",
		16#43ba# => X"b337f600",
		16#43bb# => X"33b7e600",
		16#43bc# => X"3367f700",
		16#43bd# => X"8327c102",
		16#43be# => X"232cc102",
		16#43bf# => X"330efe00",
		16#43c0# => X"3307c701",
		16#43c1# => X"232ee102",
		16#43c2# => X"13840500",
		16#43c3# => X"6ff05fb8",
		16#43c4# => X"b7860000",
		16#43c5# => X"9386f6ff",
		16#43c6# => X"e38cd5de",
		16#43c7# => X"1347f7ff",
		16#43c8# => X"93074007",
		16#43c9# => X"63d0e704",
		16#43ca# => X"232e0100",
		16#43cb# => X"232c0100",
		16#43cc# => X"232a0100",
		16#43cd# => X"93071000",
		16#43ce# => X"6f008012",
		16#43cf# => X"b7860000",
		16#43d0# => X"9386f6ff",
		16#43d1# => X"e386d5dc",
		16#43d2# => X"8327c101",
		16#43d3# => X"b7060800",
		16#43d4# => X"b3e7d700",
		16#43d5# => X"232ef100",
		16#43d6# => X"9307c0f8",
		16#43d7# => X"e346f7fc",
		16#43d8# => X"3307e040",
		16#43d9# => X"93565740",
		16#43da# => X"93080000",
		16#43db# => X"1377f701",
		16#43dc# => X"93070000",
		16#43dd# => X"13952700",
		16#43de# => X"6390d702",
		16#43df# => X"63140704",
		16#43e0# => X"93063000",
		16#43e1# => X"b386f640",
		16#43e2# => X"63d2e602",
		16#43e3# => X"13074000",
		16#43e4# => X"b307f740",
		16#43e5# => X"6f00c007",
		16#43e6# => X"3305a800",
		16#43e7# => X"03250500",
		16#43e8# => X"93871700",
		16#43e9# => X"b3e8a800",
		16#43ea# => X"6ff0dffc",
		16#43eb# => X"3303a600",
		16#43ec# => X"03230300",
		16#43ed# => X"13071700",
		16#43ee# => X"13064600",
		16#43ef# => X"232e66fe",
		16#43f0# => X"6ff09ffc",
		16#43f1# => X"93060104",
		16#43f2# => X"b386a600",
		16#43f3# => X"83a606fd",
		16#43f4# => X"130e0002",
		16#43f5# => X"330eee40",
		16#43f6# => X"b396c601",
		16#43f7# => X"b3e8d800",
		16#43f8# => X"93063000",
		16#43f9# => X"930e0000",
		16#43fa# => X"b386f640",
		16#43fb# => X"63c6de02",
		16#43fc# => X"13064000",
		16#43fd# => X"b307f640",
		16#43fe# => X"93962600",
		16#43ff# => X"13060104",
		16#4400# => X"b306d600",
		16#4401# => X"0326c101",
		16#4402# => X"3357e600",
		16#4403# => X"23a8e6fc",
		16#4404# => X"93064000",
		16#4405# => X"6f00c003",
		16#4406# => X"330fa600",
		16#4407# => X"03230f00",
		16#4408# => X"032f4f00",
		16#4409# => X"938e1e00",
		16#440a# => X"3353e300",
		16#440b# => X"331fcf01",
		16#440c# => X"3363e301",
		16#440d# => X"23206600",
		16#440e# => X"13064600",
		16#440f# => X"6ff01ffb",
		16#4410# => X"13972700",
		16#4411# => X"3307e800",
		16#4412# => X"23200700",
		16#4413# => X"93871700",
		16#4414# => X"e398d7fe",
		16#4415# => X"03270101",
		16#4416# => X"b3371001",
		16#4417# => X"b367f700",
		16#4418# => X"2328f100",
		16#4419# => X"83260102",
		16#441a# => X"83270101",
		16#441b# => X"03274102",
		16#441c# => X"03258101",
		16#441d# => X"b387f600",
		16#441e# => X"b3b6d700",
		16#441f# => X"2328f102",
		16#4420# => X"83274101",
		16#4421# => X"0328c101",
		16#4422# => X"b307f700",
		16#4423# => X"3386d700",
		16#4424# => X"33b7e700",
		16#4425# => X"b337d600",
		16#4426# => X"b367f700",
		16#4427# => X"03278102",
		16#4428# => X"8326c102",
		16#4429# => X"232ac102",
		16#442a# => X"3305a700",
		16#442b# => X"3306f500",
		16#442c# => X"3337e500",
		16#442d# => X"b337f600",
		16#442e# => X"b3860601",
		16#442f# => X"3367f700",
		16#4430# => X"232cc102",
		16#4431# => X"3387e600",
		16#4432# => X"6ff0dfe3",
		16#4433# => X"378f0000",
		16#4434# => X"13051400",
		16#4435# => X"930effff",
		16#4436# => X"b372d501",
		16#4437# => X"930f1000",
		16#4438# => X"03274102",
		16#4439# => X"03268102",
		16#443a# => X"0328c102",
		16#443b# => X"83254101",
		16#443c# => X"032e8101",
		16#443d# => X"0323c101",
		16#443e# => X"93080103",
		16#443f# => X"63c65f14",
		16#4440# => X"33e5c501",
		16#4441# => X"33656500",
		16#4442# => X"3365d500",
		16#4443# => X"6316040a",
		16#4444# => X"631c0500",
		16#4445# => X"2328f102",
		16#4446# => X"232ae102",
		16#4447# => X"232cc102",
		16#4448# => X"232e0103",
		16#4449# => X"6ff0dfc0",
		16#444a# => X"3365c700",
		16#444b# => X"33650501",
		16#444c# => X"3365f500",
		16#444d# => X"631c0500",
		16#444e# => X"2328d102",
		16#444f# => X"232ab102",
		16#4450# => X"232cc103",
		16#4451# => X"232e6102",
		16#4452# => X"6ff09fbe",
		16#4453# => X"b387f600",
		16#4454# => X"3307b700",
		16#4455# => X"2328f102",
		16#4456# => X"b3b7d700",
		16#4457# => X"b306f700",
		16#4458# => X"232ad102",
		16#4459# => X"3337b700",
		16#445a# => X"b3b6f600",
		16#445b# => X"b366d700",
		16#445c# => X"b305c601",
		16#445d# => X"b387d500",
		16#445e# => X"33b6c501",
		16#445f# => X"b3b6d700",
		16#4460# => X"b366d600",
		16#4461# => X"33066800",
		16#4462# => X"3386c600",
		16#4463# => X"232cf102",
		16#4464# => X"9317c600",
		16#4465# => X"63c60700",
		16#4466# => X"232ec102",
		16#4467# => X"6ff05fb9",
		16#4468# => X"b706f8ff",
		16#4469# => X"9386f6ff",
		16#446a# => X"3376d600",
		16#446b# => X"232ec102",
		16#446c# => X"13041000",
		16#446d# => X"6ff0dfb7",
		16#446e# => X"631e0500",
		16#446f# => X"2328f102",
		16#4470# => X"232ae102",
		16#4471# => X"232cc102",
		16#4472# => X"232e0103",
		16#4473# => X"13840e00",
		16#4474# => X"6ff01fb6",
		16#4475# => X"3366c700",
		16#4476# => X"33660601",
		16#4477# => X"b367f600",
		16#4478# => X"639c0700",
		16#4479# => X"2328d102",
		16#447a# => X"232ab102",
		16#447b# => X"232cc103",
		16#447c# => X"232e6102",
		16#447d# => X"6ff09ffd",
		16#447e# => X"232ee103",
		16#447f# => X"232c0102",
		16#4480# => X"232a0102",
		16#4481# => X"23280102",
		16#4482# => X"1307c103",
		16#4483# => X"83270700",
		16#4484# => X"8326c7ff",
		16#4485# => X"1307c7ff",
		16#4486# => X"93973700",
		16#4487# => X"93d6d601",
		16#4488# => X"b3e7d700",
		16#4489# => X"2322f700",
		16#448a# => X"e392e8fe",
		16#448b# => X"83270103",
		16#448c# => X"37840000",
		16#448d# => X"1304f4ff",
		16#448e# => X"93973700",
		16#448f# => X"2328f102",
		16#4490# => X"130a0000",
		16#4491# => X"6ff0dfae",
		16#4492# => X"b387f600",
		16#4493# => X"3307b700",
		16#4494# => X"2328f102",
		16#4495# => X"b3b7d700",
		16#4496# => X"b306f700",
		16#4497# => X"232ad102",
		16#4498# => X"3337b700",
		16#4499# => X"b3b6f600",
		16#449a# => X"b366d700",
		16#449b# => X"3306c601",
		16#449c# => X"3307d600",
		16#449d# => X"b336d700",
		16#449e# => X"3336c601",
		16#449f# => X"3366d600",
		16#44a0# => X"b3066800",
		16#44a1# => X"3306d600",
		16#44a2# => X"232ce102",
		16#44a3# => X"232ec102",
		16#44a4# => X"93870800",
		16#44a5# => X"93060000",
		16#44a6# => X"93053000",
		16#44a7# => X"03a70700",
		16#44a8# => X"03a64700",
		16#44a9# => X"93861600",
		16#44aa# => X"13571700",
		16#44ab# => X"1316f601",
		16#44ac# => X"3367c700",
		16#44ad# => X"23a0e700",
		16#44ae# => X"93874700",
		16#44af# => X"e390b6fe",
		16#44b0# => X"8327c103",
		16#44b1# => X"13040500",
		16#44b2# => X"93d71700",
		16#44b3# => X"232ef102",
		16#44b4# => X"b7870000",
		16#44b5# => X"9387f7ff",
		16#44b6# => X"e31cf4a4",
		16#44b7# => X"232e0102",
		16#44b8# => X"232c0102",
		16#44b9# => X"232a0102",
		16#44ba# => X"23280102",
		16#44bb# => X"6ff05fa4",
		16#44bc# => X"6352e028",
		16#44bd# => X"639e050c",
		16#44be# => X"03254102",
		16#44bf# => X"83258102",
		16#44c0# => X"032ec102",
		16#44c1# => X"3368b500",
		16#44c2# => X"3368c801",
		16#44c3# => X"3368f800",
		16#44c4# => X"630e08ee",
		16#44c5# => X"1306f7ff",
		16#44c6# => X"63180608",
		16#44c7# => X"83284101",
		16#44c8# => X"b387f640",
		16#44c9# => X"33b7f600",
		16#44ca# => X"3388a840",
		16#44cb# => X"33b30801",
		16#44cc# => X"3308e840",
		16#44cd# => X"2328f102",
		16#44ce# => X"232a0103",
		16#44cf# => X"13070000",
		16#44d0# => X"63f6f600",
		16#44d1# => X"33071541",
		16#44d2# => X"13371700",
		16#44d3# => X"03288101",
		16#44d4# => X"33676700",
		16#44d5# => X"b306b840",
		16#44d6# => X"3335d800",
		16#44d7# => X"b386e640",
		16#44d8# => X"232cd102",
		16#44d9# => X"63060700",
		16#44da# => X"b3850541",
		16#44db# => X"13b61500",
		16#44dc# => X"8327c101",
		16#44dd# => X"3366a600",
		16#44de# => X"13041000",
		16#44df# => X"b387c741",
		16#44e0# => X"3386c740",
		16#44e1# => X"232ec102",
		16#44e2# => X"8327c103",
		16#44e3# => X"1397c700",
		16#44e4# => X"e350079a",
		16#44e5# => X"37070800",
		16#44e6# => X"1307f7ff",
		16#44e7# => X"b3f7e700",
		16#44e8# => X"232ef102",
		16#44e9# => X"6f00c072",
		16#44ea# => X"b7870000",
		16#44eb# => X"9387f7ff",
		16#44ec# => X"630ef7e4",
		16#44ed# => X"93074007",
		16#44ee# => X"63d0c704",
		16#44ef# => X"23260102",
		16#44f0# => X"23240102",
		16#44f1# => X"23220102",
		16#44f2# => X"93071000",
		16#44f3# => X"6f008012",
		16#44f4# => X"b7870000",
		16#44f5# => X"9387f7ff",
		16#44f6# => X"6306f4f6",
		16#44f7# => X"8327c102",
		16#44f8# => X"b7060800",
		16#44f9# => X"b3e7d700",
		16#44fa# => X"2326f102",
		16#44fb# => X"93074007",
		16#44fc# => X"e3c6e7fc",
		16#44fd# => X"13060700",
		16#44fe# => X"13575640",
		16#44ff# => X"93050000",
		16#4500# => X"1376f601",
		16#4501# => X"93070000",
		16#4502# => X"93962700",
		16#4503# => X"6390e702",
		16#4504# => X"63140604",
		16#4505# => X"13073000",
		16#4506# => X"3307f740",
		16#4507# => X"6352c702",
		16#4508# => X"13074000",
		16#4509# => X"b307f740",
		16#450a# => X"6f00c007",
		16#450b# => X"b386d800",
		16#450c# => X"83a60600",
		16#450d# => X"93871700",
		16#450e# => X"b3e5d500",
		16#450f# => X"6ff0dffc",
		16#4510# => X"3305d300",
		16#4511# => X"03250500",
		16#4512# => X"13061600",
		16#4513# => X"13034300",
		16#4514# => X"232ea3fe",
		16#4515# => X"6ff09ffc",
		16#4516# => X"13070104",
		16#4517# => X"3307d700",
		16#4518# => X"032707fe",
		16#4519# => X"13080002",
		16#451a# => X"3308c840",
		16#451b# => X"33170701",
		16#451c# => X"b3e5e500",
		16#451d# => X"13073000",
		16#451e# => X"130e0000",
		16#451f# => X"3307f740",
		16#4520# => X"6346ee02",
		16#4521# => X"93064000",
		16#4522# => X"b387f640",
		16#4523# => X"13172700",
		16#4524# => X"93060104",
		16#4525# => X"3387e600",
		16#4526# => X"8326c102",
		16#4527# => X"33d6c600",
		16#4528# => X"2320c7fe",
		16#4529# => X"93064000",
		16#452a# => X"6f00c003",
		16#452b# => X"b30ed300",
		16#452c# => X"03a50e00",
		16#452d# => X"83ae4e00",
		16#452e# => X"130e1e00",
		16#452f# => X"3355c500",
		16#4530# => X"b39e0e01",
		16#4531# => X"3365d501",
		16#4532# => X"2320a300",
		16#4533# => X"13034300",
		16#4534# => X"6ff01ffb",
		16#4535# => X"13972700",
		16#4536# => X"3387e800",
		16#4537# => X"23200700",
		16#4538# => X"93871700",
		16#4539# => X"e398d7fe",
		16#453a# => X"03270102",
		16#453b# => X"b337b000",
		16#453c# => X"b367f700",
		16#453d# => X"2320f102",
		16#453e# => X"83264101",
		16#453f# => X"83250101",
		16#4540# => X"03270102",
		16#4541# => X"83274102",
		16#4542# => X"3387e540",
		16#4543# => X"b387f640",
		16#4544# => X"33b6f600",
		16#4545# => X"b3b6e500",
		16#4546# => X"b386d740",
		16#4547# => X"232ad102",
		16#4548# => X"2328e102",
		16#4549# => X"93060000",
		16#454a# => X"63f4e500",
		16#454b# => X"93b61700",
		16#454c# => X"b3e6c600",
		16#454d# => X"03278102",
		16#454e# => X"03268101",
		16#454f# => X"3307e640",
		16#4550# => X"b307d740",
		16#4551# => X"232cf102",
		16#4552# => X"b335e600",
		16#4553# => X"13060000",
		16#4554# => X"63840600",
		16#4555# => X"13361700",
		16#4556# => X"8327c101",
		16#4557# => X"0327c102",
		16#4558# => X"3366b600",
		16#4559# => X"b387e740",
		16#455a# => X"b387c740",
		16#455b# => X"232ef102",
		16#455c# => X"6ff09fe1",
		16#455d# => X"630c0728",
		16#455e# => X"631a040e",
		16#455f# => X"03234101",
		16#4560# => X"83288101",
		16#4561# => X"832ec101",
		16#4562# => X"336e1301",
		16#4563# => X"336ede01",
		16#4564# => X"336ede00",
		16#4565# => X"63160e02",
		16#4566# => X"2328f102",
		16#4567# => X"83274102",
		16#4568# => X"13840500",
		16#4569# => X"232af102",
		16#456a# => X"83278102",
		16#456b# => X"232cf102",
		16#456c# => X"8327c102",
		16#456d# => X"232ef102",
		16#456e# => X"130a0500",
		16#456f# => X"6ff04ff7",
		16#4570# => X"130ef0ff",
		16#4571# => X"631ec707",
		16#4572# => X"03284102",
		16#4573# => X"b386d740",
		16#4574# => X"33b7d700",
		16#4575# => X"33066840",
		16#4576# => X"333ec800",
		16#4577# => X"3306e640",
		16#4578# => X"2328d102",
		16#4579# => X"232ac102",
		16#457a# => X"13070000",
		16#457b# => X"63f6d700",
		16#457c# => X"33070341",
		16#457d# => X"13371700",
		16#457e# => X"03288102",
		16#457f# => X"3367c701",
		16#4580# => X"93060000",
		16#4581# => X"33061841",
		16#4582# => X"3333c800",
		16#4583# => X"3306e640",
		16#4584# => X"232cc102",
		16#4585# => X"63060700",
		16#4586# => X"b3880841",
		16#4587# => X"93b61800",
		16#4588# => X"8327c102",
		16#4589# => X"b3e86600",
		16#458a# => X"b387d741",
		16#458b# => X"b3871741",
		16#458c# => X"232ef102",
		16#458d# => X"13840500",
		16#458e# => X"130a0500",
		16#458f# => X"6ff0dfd4",
		16#4590# => X"b7860000",
		16#4591# => X"9386f6ff",
		16#4592# => X"e388d5f4",
		16#4593# => X"1347f7ff",
		16#4594# => X"93074007",
		16#4595# => X"63d0e704",
		16#4596# => X"232e0100",
		16#4597# => X"232c0100",
		16#4598# => X"232a0100",
		16#4599# => X"93071000",
		16#459a# => X"6f008012",
		16#459b# => X"b7860000",
		16#459c# => X"9386f6ff",
		16#459d# => X"e382d5f2",
		16#459e# => X"8327c101",
		16#459f# => X"b7060800",
		16#45a0# => X"b3e7d700",
		16#45a1# => X"232ef100",
		16#45a2# => X"9307c0f8",
		16#45a3# => X"e346f7fc",
		16#45a4# => X"3307e040",
		16#45a5# => X"93565740",
		16#45a6# => X"13030000",
		16#45a7# => X"1377f701",
		16#45a8# => X"93070000",
		16#45a9# => X"93982700",
		16#45aa# => X"6390d702",
		16#45ab# => X"63140704",
		16#45ac# => X"93063000",
		16#45ad# => X"b386f640",
		16#45ae# => X"63d2e602",
		16#45af# => X"13074000",
		16#45b0# => X"b307f740",
		16#45b1# => X"6f00c007",
		16#45b2# => X"b3081801",
		16#45b3# => X"83a80800",
		16#45b4# => X"93871700",
		16#45b5# => X"33631301",
		16#45b6# => X"6ff0dffc",
		16#45b7# => X"330e1601",
		16#45b8# => X"032e0e00",
		16#45b9# => X"13071700",
		16#45ba# => X"13064600",
		16#45bb# => X"232ec6ff",
		16#45bc# => X"6ff09ffc",
		16#45bd# => X"93060104",
		16#45be# => X"b3861601",
		16#45bf# => X"83a606fd",
		16#45c0# => X"930e0002",
		16#45c1# => X"b38eee40",
		16#45c2# => X"b396d601",
		16#45c3# => X"3363d300",
		16#45c4# => X"93063000",
		16#45c5# => X"130f0000",
		16#45c6# => X"b386f640",
		16#45c7# => X"6346df02",
		16#45c8# => X"13064000",
		16#45c9# => X"b307f640",
		16#45ca# => X"93962600",
		16#45cb# => X"13060104",
		16#45cc# => X"b306d600",
		16#45cd# => X"0326c101",
		16#45ce# => X"3357e600",
		16#45cf# => X"23a8e6fc",
		16#45d0# => X"93064000",
		16#45d1# => X"6f00c003",
		16#45d2# => X"b30f1601",
		16#45d3# => X"03ae0f00",
		16#45d4# => X"83af4f00",
		16#45d5# => X"130f1f00",
		16#45d6# => X"335eee00",
		16#45d7# => X"b39fdf01",
		16#45d8# => X"336efe01",
		16#45d9# => X"2320c601",
		16#45da# => X"13064600",
		16#45db# => X"6ff01ffb",
		16#45dc# => X"13972700",
		16#45dd# => X"3307e800",
		16#45de# => X"23200700",
		16#45df# => X"93871700",
		16#45e0# => X"e398d7fe",
		16#45e1# => X"03270101",
		16#45e2# => X"b3376000",
		16#45e3# => X"b367f700",
		16#45e4# => X"2328f100",
		16#45e5# => X"83264102",
		16#45e6# => X"03280102",
		16#45e7# => X"03270101",
		16#45e8# => X"83274101",
		16#45e9# => X"3307e840",
		16#45ea# => X"b387f640",
		16#45eb# => X"33b6f600",
		16#45ec# => X"b336e800",
		16#45ed# => X"b386d740",
		16#45ee# => X"232ad102",
		16#45ef# => X"2328e102",
		16#45f0# => X"93060000",
		16#45f1# => X"6374e800",
		16#45f2# => X"93b61700",
		16#45f3# => X"b3e6c600",
		16#45f4# => X"03278101",
		16#45f5# => X"03268102",
		16#45f6# => X"3307e640",
		16#45f7# => X"b307d740",
		16#45f8# => X"232cf102",
		16#45f9# => X"3338e600",
		16#45fa# => X"13060000",
		16#45fb# => X"63840600",
		16#45fc# => X"13361700",
		16#45fd# => X"8327c102",
		16#45fe# => X"0327c101",
		16#45ff# => X"33660601",
		16#4600# => X"b387e740",
		16#4601# => X"b387c740",
		16#4602# => X"6ff09fe2",
		16#4603# => X"b78f0000",
		16#4604# => X"930e1400",
		16#4605# => X"9382ffff",
		16#4606# => X"b3fe5e00",
		16#4607# => X"130f1000",
		16#4608# => X"83254102",
		16#4609# => X"03264101",
		16#460a# => X"03288101",
		16#460b# => X"032ec101",
		16#460c# => X"83288102",
		16#460d# => X"0323c102",
		16#460e# => X"634edf1d",
		16#460f# => X"b3ee1501",
		16#4610# => X"336f0601",
		16#4611# => X"b3ee6e00",
		16#4612# => X"336fcf01",
		16#4613# => X"b3eefe00",
		16#4614# => X"336fdf00",
		16#4615# => X"63180410",
		16#4616# => X"63120f02",
		16#4617# => X"2328f102",
		16#4618# => X"232ab102",
		16#4619# => X"232c1103",
		16#461a# => X"232e6102",
		16#461b# => X"e3960ed4",
		16#461c# => X"13040000",
		16#461d# => X"130a0000",
		16#461e# => X"6ff08fd0",
		16#461f# => X"639c0e00",
		16#4620# => X"2328d102",
		16#4621# => X"232ac102",
		16#4622# => X"232c0103",
		16#4623# => X"232ec103",
		16#4624# => X"6ff00fca",
		16#4625# => X"b38ef640",
		16#4626# => X"b302b640",
		16#4627# => X"b3bfd601",
		16#4628# => X"333f5600",
		16#4629# => X"b382f241",
		16#462a# => X"2328d103",
		16#462b# => X"232a5102",
		16#462c# => X"930f0000",
		16#462d# => X"63f6d601",
		16#462e# => X"b38fc540",
		16#462f# => X"93bf1f00",
		16#4630# => X"b3031841",
		16#4631# => X"b3efef01",
		16#4632# => X"b389f341",
		16#4633# => X"232c3103",
		16#4634# => X"b33a7800",
		16#4635# => X"13090000",
		16#4636# => X"63840f00",
		16#4637# => X"13b91300",
		16#4638# => X"330f6e40",
		16#4639# => X"33695901",
		16#463a# => X"330f2f41",
		16#463b# => X"232ee103",
		16#463c# => X"931fcf00",
		16#463d# => X"63de0f04",
		16#463e# => X"b386d740",
		16#463f# => X"3386c540",
		16#4640# => X"b3bed700",
		16#4641# => X"b30ed641",
		16#4642# => X"232ad103",
		16#4643# => X"2328d102",
		16#4644# => X"b3b5c500",
		16#4645# => X"930e0000",
		16#4646# => X"63f4d700",
		16#4647# => X"933e1600",
		16#4648# => X"b3870841",
		16#4649# => X"b3e5be00",
		16#464a# => X"b3b6f800",
		16#464b# => X"b387b740",
		16#464c# => X"232cf102",
		16#464d# => X"63840500",
		16#464e# => X"13b71300",
		16#464f# => X"3303c341",
		16#4650# => X"3367d700",
		16#4651# => X"3303e340",
		16#4652# => X"232e6102",
		16#4653# => X"6ff0dfc6",
		16#4654# => X"b3ee5e00",
		16#4655# => X"b3ee3e01",
		16#4656# => X"b3eeee01",
		16#4657# => X"e38a0ef0",
		16#4658# => X"6ff00fbd",
		16#4659# => X"93030103",
		16#465a# => X"631e0f04",
		16#465b# => X"639e0e02",
		16#465c# => X"232ef103",
		16#465d# => X"232c0102",
		16#465e# => X"232a0102",
		16#465f# => X"23280102",
		16#4660# => X"9307c103",
		16#4661# => X"03a70700",
		16#4662# => X"83a6c7ff",
		16#4663# => X"9387c7ff",
		16#4664# => X"13173700",
		16#4665# => X"93d6d601",
		16#4666# => X"3367d700",
		16#4667# => X"23a2e700",
		16#4668# => X"e392f3fe",
		16#4669# => X"6ff09f88",
		16#466a# => X"2328f102",
		16#466b# => X"232ab102",
		16#466c# => X"232c1103",
		16#466d# => X"232e6102",
		16#466e# => X"130a0500",
		16#466f# => X"13840200",
		16#4670# => X"6ff00fb7",
		16#4671# => X"639c0e00",
		16#4672# => X"2328d102",
		16#4673# => X"232ac102",
		16#4674# => X"232c0103",
		16#4675# => X"232ec103",
		16#4676# => X"6ff05ffe",
		16#4677# => X"232ef103",
		16#4678# => X"232c0102",
		16#4679# => X"232a0102",
		16#467a# => X"23280102",
		16#467b# => X"9307c103",
		16#467c# => X"03a70700",
		16#467d# => X"83a6c7ff",
		16#467e# => X"9387c7ff",
		16#467f# => X"13173700",
		16#4680# => X"93d6d601",
		16#4681# => X"3367d700",
		16#4682# => X"23a2e700",
		16#4683# => X"e392f3fe",
		16#4684# => X"6ff0df81",
		16#4685# => X"b38ef640",
		16#4686# => X"b302b640",
		16#4687# => X"b3bfd601",
		16#4688# => X"333f5600",
		16#4689# => X"b382f241",
		16#468a# => X"2328d103",
		16#468b# => X"232a5102",
		16#468c# => X"930f0000",
		16#468d# => X"63f6d601",
		16#468e# => X"b38fc540",
		16#468f# => X"93bf1f00",
		16#4690# => X"b3031841",
		16#4691# => X"b3efef01",
		16#4692# => X"b389f341",
		16#4693# => X"232c3103",
		16#4694# => X"b33a7800",
		16#4695# => X"13090000",
		16#4696# => X"63840f00",
		16#4697# => X"13b91300",
		16#4698# => X"330f6e40",
		16#4699# => X"33695901",
		16#469a# => X"330f2f41",
		16#469b# => X"232ee103",
		16#469c# => X"931fcf00",
		16#469d# => X"63d00f0e",
		16#469e# => X"b386d740",
		16#469f# => X"3386c540",
		16#46a0# => X"b3bed700",
		16#46a1# => X"b30ed641",
		16#46a2# => X"232ad103",
		16#46a3# => X"2328d102",
		16#46a4# => X"b3b5c500",
		16#46a5# => X"930e0000",
		16#46a6# => X"63f4d700",
		16#46a7# => X"933e1600",
		16#46a8# => X"b3870841",
		16#46a9# => X"b3e5be00",
		16#46aa# => X"b3b6f800",
		16#46ab# => X"b387b740",
		16#46ac# => X"232cf102",
		16#46ad# => X"63840500",
		16#46ae# => X"13b71300",
		16#46af# => X"3303c341",
		16#46b0# => X"3367d700",
		16#46b1# => X"3307e340",
		16#46b2# => X"232ee102",
		16#46b3# => X"130a0500",
		16#46b4# => X"0325c103",
		16#46b5# => X"630a0508",
		16#46b6# => X"ef001043",
		16#46b7# => X"930a45ff",
		16#46b8# => X"13d9fa41",
		16#46b9# => X"b7090080",
		16#46ba# => X"1379f901",
		16#46bb# => X"9389f901",
		16#46bc# => X"33095901",
		16#46bd# => X"b3f93a01",
		16#46be# => X"13595940",
		16#46bf# => X"63d80900",
		16#46c0# => X"9389f9ff",
		16#46c1# => X"93e909fe",
		16#46c2# => X"93891900",
		16#46c3# => X"638a0908",
		16#46c4# => X"9305c0ff",
		16#46c5# => X"13050900",
		16#46c6# => X"ef009031",
		16#46c7# => X"93060002",
		16#46c8# => X"13172900",
		16#46c9# => X"130800ff",
		16#46ca# => X"b3863641",
		16#46cb# => X"1305c5ff",
		16#46cc# => X"6312050b",
		16#46cd# => X"93070104",
		16#46ce# => X"3387e700",
		16#46cf# => X"83270103",
		16#46d0# => X"1309f9ff",
		16#46d1# => X"b3993701",
		16#46d2# => X"232837ff",
		16#46d3# => X"1307f0ff",
		16#46d4# => X"6f00400c",
		16#46d5# => X"b3ee5e00",
		16#46d6# => X"b3ee3e01",
		16#46d7# => X"b3eeee01",
		16#46d8# => X"e3880ed0",
		16#46d9# => X"6ff0dff6",
		16#46da# => X"03258103",
		16#46db# => X"63080500",
		16#46dc# => X"ef009039",
		16#46dd# => X"13050502",
		16#46de# => X"6ff05ff6",
		16#46df# => X"03254103",
		16#46e0# => X"63080500",
		16#46e1# => X"ef005038",
		16#46e2# => X"13050504",
		16#46e3# => X"6ff01ff5",
		16#46e4# => X"03250103",
		16#46e5# => X"ef005037",
		16#46e6# => X"13050506",
		16#46e7# => X"6ff01ff4",
		16#46e8# => X"9305c0ff",
		16#46e9# => X"13050900",
		16#46ea# => X"ef009028",
		16#46eb# => X"93090103",
		16#46ec# => X"93073000",
		16#46ed# => X"3387a900",
		16#46ee# => X"0327c700",
		16#46ef# => X"9387f7ff",
		16#46f0# => X"9389c9ff",
		16#46f1# => X"23a8e900",
		16#46f2# => X"e3d627ff",
		16#46f3# => X"1309f9ff",
		16#46f4# => X"6ff0dff7",
		16#46f5# => X"93070103",
		16#46f6# => X"b385a700",
		16#46f7# => X"3306a700",
		16#46f8# => X"3386c700",
		16#46f9# => X"83a7c500",
		16#46fa# => X"83a50501",
		16#46fb# => X"b3d7d700",
		16#46fc# => X"b3953501",
		16#46fd# => X"b3e7b700",
		16#46fe# => X"2328f600",
		16#46ff# => X"6ff01ff3",
		16#4700# => X"93172900",
		16#4701# => X"93060103",
		16#4702# => X"b387f600",
		16#4703# => X"23a00700",
		16#4704# => X"1309f9ff",
		16#4705# => X"e316e9fe",
		16#4706# => X"63c08a16",
		16#4707# => X"33848a40",
		16#4708# => X"13041400",
		16#4709# => X"9357f441",
		16#470a# => X"37070080",
		16#470b# => X"93f7f701",
		16#470c# => X"1307f701",
		16#470d# => X"b3878700",
		16#470e# => X"3374e400",
		16#470f# => X"93d75740",
		16#4710# => X"63580400",
		16#4711# => X"1304f4ff",
		16#4712# => X"136404fe",
		16#4713# => X"13041400",
		16#4714# => X"93060400",
		16#4715# => X"13050000",
		16#4716# => X"13070000",
		16#4717# => X"634af702",
		16#4718# => X"13870700",
		16#4719# => X"63d40700",
		16#471a# => X"13070000",
		16#471b# => X"13932700",
		16#471c# => X"631a0404",
		16#471d# => X"13063000",
		16#471e# => X"13070103",
		16#471f# => X"3306f640",
		16#4720# => X"6356d602",
		16#4721# => X"13074000",
		16#4722# => X"b307f740",
		16#4723# => X"6f00c008",
		16#4724# => X"13162700",
		16#4725# => X"93050103",
		16#4726# => X"3386c500",
		16#4727# => X"03260600",
		16#4728# => X"13071700",
		16#4729# => X"3365c500",
		16#472a# => X"6ff05ffb",
		16#472b# => X"b3056700",
		16#472c# => X"83a50500",
		16#472d# => X"93861600",
		16#472e# => X"13074700",
		16#472f# => X"232eb7fe",
		16#4730# => X"6ff01ffc",
		16#4731# => X"13172700",
		16#4732# => X"93060104",
		16#4733# => X"3387e600",
		16#4734# => X"032707ff",
		16#4735# => X"13060002",
		16#4736# => X"33068640",
		16#4737# => X"3317c700",
		16#4738# => X"3365e500",
		16#4739# => X"13073000",
		16#473a# => X"93050103",
		16#473b# => X"13080000",
		16#473c# => X"3307f740",
		16#473d# => X"6346e802",
		16#473e# => X"93064000",
		16#473f# => X"b387f640",
		16#4740# => X"13172700",
		16#4741# => X"93060104",
		16#4742# => X"3387e600",
		16#4743# => X"8326c103",
		16#4744# => X"33d48600",
		16#4745# => X"232887fe",
		16#4746# => X"93063000",
		16#4747# => X"6f000004",
		16#4748# => X"b3886500",
		16#4749# => X"83a60800",
		16#474a# => X"83a84800",
		16#474b# => X"13081800",
		16#474c# => X"b3d68600",
		16#474d# => X"b398c800",
		16#474e# => X"b3e61601",
		16#474f# => X"23a0d500",
		16#4750# => X"93854500",
		16#4751# => X"6ff01ffb",
		16#4752# => X"13972700",
		16#4753# => X"13060103",
		16#4754# => X"3307e600",
		16#4755# => X"23200700",
		16#4756# => X"93871700",
		16#4757# => X"e3d6f6fe",
		16#4758# => X"03270103",
		16#4759# => X"b337a000",
		16#475a# => X"13040000",
		16#475b# => X"b367f700",
		16#475c# => X"2328f102",
		16#475d# => X"6fe0dffb",
		16#475e# => X"8327c103",
		16#475f# => X"3707f8ff",
		16#4760# => X"1307f7ff",
		16#4761# => X"33045441",
		16#4762# => X"b3f7e700",
		16#4763# => X"6fe01fdd",
		16#4764# => X"232e0102",
		16#4765# => X"232c0102",
		16#4766# => X"232a0102",
		16#4767# => X"23280102",
		16#4768# => X"6ff00f81",
		16#4769# => X"03274500",
		16#476a# => X"83278500",
		16#476b# => X"0326c500",
		16#476c# => X"83260500",
		16#476d# => X"130101fe",
		16#476e# => X"2322e100",
		16#476f# => X"2324f100",
		16#4770# => X"232ae100",
		16#4771# => X"232cf100",
		16#4772# => X"37470000",
		16#4773# => X"93171600",
		16#4774# => X"2320d100",
		16#4775# => X"2328d100",
		16#4776# => X"2326c100",
		16#4777# => X"93d61701",
		16#4778# => X"9307e7ff",
		16#4779# => X"13050000",
		16#477a# => X"63d0d702",
		16#477b# => X"9307d701",
		16#477c# => X"93150601",
		16#477d# => X"1356f601",
		16#477e# => X"63dcd700",
		16#477f# => X"37050080",
		16#4780# => X"1345f5ff",
		16#4781# => X"3305a600",
		16#4782# => X"13010102",
		16#4783# => X"67800000",
		16#4784# => X"b7070100",
		16#4785# => X"93d50501",
		16#4786# => X"b3e5f500",
		16#4787# => X"9307f706",
		16#4788# => X"b387d740",
		16#4789# => X"13d75740",
		16#478a# => X"232eb100",
		16#478b# => X"93f7f701",
		16#478c# => X"6392070a",
		16#478d# => X"93053000",
		16#478e# => X"93060101",
		16#478f# => X"13152700",
		16#4790# => X"b385e540",
		16#4791# => X"63def502",
		16#4792# => X"93074000",
		16#4793# => X"3387e740",
		16#4794# => X"93060101",
		16#4795# => X"93172700",
		16#4796# => X"b387f600",
		16#4797# => X"93064000",
		16#4798# => X"23a00700",
		16#4799# => X"13071700",
		16#479a# => X"93874700",
		16#479b# => X"e31ad7fe",
		16#479c# => X"03250101",
		16#479d# => X"e30a06f8",
		16#479e# => X"3305a040",
		16#479f# => X"6ff0dff8",
		16#47a0# => X"3388a600",
		16#47a1# => X"03280800",
		16#47a2# => X"93871700",
		16#47a3# => X"93864600",
		16#47a4# => X"23ae06ff",
		16#47a5# => X"6ff01ffb",
		16#47a6# => X"832605ff",
		16#47a7# => X"032307ff",
		16#47a8# => X"b3961601",
		16#47a9# => X"3353f300",
		16#47aa# => X"b3e66600",
		16#47ab# => X"2328d100",
		16#47ac# => X"93061000",
		16#47ad# => X"e3c206ff",
		16#47ae# => X"13871600",
		16#47af# => X"13050102",
		16#47b0# => X"93962600",
		16#47b1# => X"b306d500",
		16#47b2# => X"b3d7f500",
		16#47b3# => X"23a8f6fe",
		16#47b4# => X"6ff01ff8",
		16#47b5# => X"13051700",
		16#47b6# => X"93080102",
		16#47b7# => X"13083000",
		16#47b8# => X"13152500",
		16#47b9# => X"3308e840",
		16#47ba# => X"3385a800",
		16#47bb# => X"13172700",
		16#47bc# => X"93080002",
		16#47bd# => X"13030102",
		16#47be# => X"93060000",
		16#47bf# => X"b388f840",
		16#47c0# => X"3307e300",
		16#47c1# => X"6ff01ffb",
		16#47c2# => X"130101fd",
		16#47c3# => X"23229102",
		16#47c4# => X"23261102",
		16#47c5# => X"23248102",
		16#47c6# => X"23202103",
		16#47c7# => X"93040500",
		16#47c8# => X"63860514",
		16#47c9# => X"13840500",
		16#47ca# => X"13d9f501",
		16#47cb# => X"63d40500",
		16#47cc# => X"3304b040",
		16#47cd# => X"13050400",
		16#47ce# => X"ef00007d",
		16#47cf# => X"93051505",
		16#47d0# => X"b7470000",
		16#47d1# => X"9387e701",
		16#47d2# => X"13d75540",
		16#47d3# => X"23288100",
		16#47d4# => X"232a0100",
		16#47d5# => X"232c0100",
		16#47d6# => X"232e0100",
		16#47d7# => X"93f5f501",
		16#47d8# => X"b387a740",
		16#47d9# => X"638c0502",
		16#47da# => X"93062000",
		16#47db# => X"631cd70e",
		16#47dc# => X"93060002",
		16#47dd# => X"b386b640",
		16#47de# => X"b356d400",
		16#47df# => X"232ed100",
		16#47e0# => X"9306f7ff",
		16#47e1# => X"13060102",
		16#47e2# => X"13172700",
		16#47e3# => X"3307e600",
		16#47e4# => X"3314b400",
		16#47e5# => X"232887fe",
		16#47e6# => X"6f004003",
		16#47e7# => X"93063000",
		16#47e8# => X"b386e640",
		16#47e9# => X"13060102",
		16#47ea# => X"93962600",
		16#47eb# => X"b306d600",
		16#47ec# => X"83a606ff",
		16#47ed# => X"13062000",
		16#47ee# => X"232ed100",
		16#47ef# => X"93062000",
		16#47f0# => X"6316c700",
		16#47f1# => X"232c8100",
		16#47f2# => X"93061000",
		16#47f3# => X"13060101",
		16#47f4# => X"13972600",
		16#47f5# => X"3307e600",
		16#47f6# => X"1306f0ff",
		16#47f7# => X"23200700",
		16#47f8# => X"9386f6ff",
		16#47f9# => X"1307c7ff",
		16#47fa# => X"e39ac6fe",
		16#47fb# => X"0327c101",
		16#47fc# => X"b7060180",
		16#47fd# => X"9386f6ff",
		16#47fe# => X"2316e100",
		16#47ff# => X"37870000",
		16#4800# => X"1307f7ff",
		16#4801# => X"b3f7e700",
		16#4802# => X"13970701",
		16#4803# => X"8327c100",
		16#4804# => X"1319f901",
		16#4805# => X"8320c102",
		16#4806# => X"b3f7d700",
		16#4807# => X"b3e7e700",
		16#4808# => X"37070080",
		16#4809# => X"1347f7ff",
		16#480a# => X"b3f7e700",
		16#480b# => X"03270101",
		16#480c# => X"03248102",
		16#480d# => X"b3e72701",
		16#480e# => X"23a0e400",
		16#480f# => X"03274101",
		16#4810# => X"23a6f400",
		16#4811# => X"13850400",
		16#4812# => X"23a2e400",
		16#4813# => X"03278101",
		16#4814# => X"03290102",
		16#4815# => X"23a4e400",
		16#4816# => X"83244102",
		16#4817# => X"13010103",
		16#4818# => X"67800000",
		16#4819# => X"13073000",
		16#481a# => X"6ff09ff1",
		16#481b# => X"232e0100",
		16#481c# => X"232c0100",
		16#481d# => X"232a0100",
		16#481e# => X"23280100",
		16#481f# => X"93070000",
		16#4820# => X"13090000",
		16#4821# => X"6ff09ff6",
		16#4822# => X"93574601",
		16#4823# => X"37071000",
		16#4824# => X"1307f7ff",
		16#4825# => X"93f7f77f",
		16#4826# => X"130101fc",
		16#4827# => X"3377c700",
		16#4828# => X"93861700",
		16#4829# => X"232c8102",
		16#482a# => X"232a9102",
		16#482b# => X"232e1102",
		16#482c# => X"9354f601",
		16#482d# => X"23282103",
		16#482e# => X"23263103",
		16#482f# => X"23244103",
		16#4830# => X"23225103",
		16#4831# => X"2328b100",
		16#4832# => X"232ae100",
		16#4833# => X"232e0100",
		16#4834# => X"232c0100",
		16#4835# => X"93f6f67f",
		16#4836# => X"13061000",
		16#4837# => X"13040500",
		16#4838# => X"635cd60a",
		16#4839# => X"b7460000",
		16#483a# => X"938606c0",
		16#483b# => X"13d54500",
		16#483c# => X"b387d700",
		16#483d# => X"93564700",
		16#483e# => X"1317c701",
		16#483f# => X"3367a700",
		16#4840# => X"9395c501",
		16#4841# => X"232ed100",
		16#4842# => X"232ce100",
		16#4843# => X"232ab100",
		16#4844# => X"23280100",
		16#4845# => X"0327c101",
		16#4846# => X"b7060180",
		16#4847# => X"9386f6ff",
		16#4848# => X"2316e100",
		16#4849# => X"37870000",
		16#484a# => X"1307f7ff",
		16#484b# => X"b3f7e700",
		16#484c# => X"0327c100",
		16#484d# => X"93970701",
		16#484e# => X"9394f401",
		16#484f# => X"3377d700",
		16#4850# => X"b367f700",
		16#4851# => X"37070080",
		16#4852# => X"1347f7ff",
		16#4853# => X"b3f7e700",
		16#4854# => X"b3e49700",
		16#4855# => X"83270101",
		16#4856# => X"23269400",
		16#4857# => X"13050400",
		16#4858# => X"2320f400",
		16#4859# => X"83274101",
		16#485a# => X"8320c103",
		16#485b# => X"83244103",
		16#485c# => X"2322f400",
		16#485d# => X"83278101",
		16#485e# => X"03290103",
		16#485f# => X"8329c102",
		16#4860# => X"2324f400",
		16#4861# => X"03248103",
		16#4862# => X"032a8102",
		16#4863# => X"832a4102",
		16#4864# => X"13010104",
		16#4865# => X"67800000",
		16#4866# => X"3365b700",
		16#4867# => X"63900710",
		16#4868# => X"e30a05f6",
		16#4869# => X"63040706",
		16#486a# => X"13050700",
		16#486b# => X"ef00c055",
		16#486c# => X"130a0500",
		16#486d# => X"93091a03",
		16#486e# => X"13d95940",
		16#486f# => X"93f9f901",
		16#4870# => X"638c0904",
		16#4871# => X"9305c0ff",
		16#4872# => X"13050900",
		16#4873# => X"ef004046",
		16#4874# => X"93070002",
		16#4875# => X"930a0101",
		16#4876# => X"130600ff",
		16#4877# => X"b3873741",
		16#4878# => X"1305c5ff",
		16#4879# => X"938acaff",
		16#487a# => X"6318c508",
		16#487b# => X"93070102",
		16#487c# => X"9306f9ff",
		16#487d# => X"13192900",
		16#487e# => X"33892701",
		16#487f# => X"83270101",
		16#4880# => X"b3993701",
		16#4881# => X"232839ff",
		16#4882# => X"6f000004",
		16#4883# => X"ef00c04f",
		16#4884# => X"130a0502",
		16#4885# => X"6ff01ffa",
		16#4886# => X"9305c0ff",
		16#4887# => X"13050900",
		16#4888# => X"ef000041",
		16#4889# => X"93090101",
		16#488a# => X"93073000",
		16#488b# => X"3387a900",
		16#488c# => X"0327c700",
		16#488d# => X"9387f7ff",
		16#488e# => X"9389c9ff",
		16#488f# => X"23a8e900",
		16#4890# => X"e3d627ff",
		16#4891# => X"9306f9ff",
		16#4892# => X"93070101",
		16#4893# => X"13972600",
		16#4894# => X"3387e700",
		16#4895# => X"9307f0ff",
		16#4896# => X"23200700",
		16#4897# => X"9386f6ff",
		16#4898# => X"1307c7ff",
		16#4899# => X"e39af6fe",
		16#489a# => X"b7470000",
		16#489b# => X"9387c7c0",
		16#489c# => X"b3874741",
		16#489d# => X"6ff01fea",
		16#489e# => X"13070101",
		16#489f# => X"b306a700",
		16#48a0# => X"03a7c600",
		16#48a1# => X"83a60601",
		16#48a2# => X"3357f700",
		16#48a3# => X"b3963601",
		16#48a4# => X"3367d700",
		16#48a5# => X"23a8ea00",
		16#48a6# => X"6ff09ff4",
		16#48a7# => X"b7870000",
		16#48a8# => X"63080502",
		16#48a9# => X"9317c701",
		16#48aa# => X"93d64500",
		16#48ab# => X"b3e7d700",
		16#48ac# => X"232cf100",
		16#48ad# => X"13574700",
		16#48ae# => X"b7870000",
		16#48af# => X"9395c501",
		16#48b0# => X"3367f700",
		16#48b1# => X"232ab100",
		16#48b2# => X"23280100",
		16#48b3# => X"232ee100",
		16#48b4# => X"9387f7ff",
		16#48b5# => X"6ff01fe4",
		16#48b6# => X"8325c500",
		16#48b7# => X"83278500",
		16#48b8# => X"03274500",
		16#48b9# => X"130101fe",
		16#48ba# => X"83260500",
		16#48bb# => X"2324f100",
		16#48bc# => X"232cf100",
		16#48bd# => X"93970501",
		16#48be# => X"2322e100",
		16#48bf# => X"232ae100",
		16#48c0# => X"93d70701",
		16#48c1# => X"13971500",
		16#48c2# => X"2326b100",
		16#48c3# => X"2320d100",
		16#48c4# => X"2328d100",
		16#48c5# => X"232ef100",
		16#48c6# => X"13571701",
		16#48c7# => X"93d5f501",
		16#48c8# => X"13030101",
		16#48c9# => X"1306c101",
		16#48ca# => X"83270600",
		16#48cb# => X"8326c6ff",
		16#48cc# => X"1306c6ff",
		16#48cd# => X"93973700",
		16#48ce# => X"93d6d601",
		16#48cf# => X"b3e7d700",
		16#48d0# => X"2322f600",
		16#48d1# => X"e312c3fe",
		16#48d2# => X"83260101",
		16#48d3# => X"93071700",
		16#48d4# => X"13953600",
		16#48d5# => X"b7860000",
		16#48d6# => X"9386f6ff",
		16#48d7# => X"b3f7d700",
		16#48d8# => X"2328a100",
		16#48d9# => X"93061000",
		16#48da# => X"63dcf61a",
		16#48db# => X"b7c7ffff",
		16#48dc# => X"93870740",
		16#48dd# => X"3307f700",
		16#48de# => X"9307e07f",
		16#48df# => X"63cee71e",
		16#48e0# => X"6358e006",
		16#48e1# => X"03288101",
		16#48e2# => X"0326c101",
		16#48e3# => X"83274101",
		16#48e4# => X"9356c801",
		16#48e5# => X"13164600",
		16#48e6# => X"3366d600",
		16#48e7# => X"93964700",
		16#48e8# => X"b3e6a600",
		16#48e9# => X"93d7c701",
		16#48ea# => X"13184800",
		16#48eb# => X"b336d000",
		16#48ec# => X"b3e70701",
		16#48ed# => X"b3e6f600",
		16#48ee# => X"232ac100",
		16#48ef# => X"2328d100",
		16#48f0# => X"83260101",
		16#48f1# => X"83274101",
		16#48f2# => X"13f67600",
		16#48f3# => X"630c061a",
		16#48f4# => X"13f6f600",
		16#48f5# => X"13054000",
		16#48f6# => X"6306a61a",
		16#48f7# => X"13864600",
		16#48f8# => X"b336d600",
		16#48f9# => X"b387d700",
		16#48fa# => X"93060600",
		16#48fb# => X"6f008019",
		16#48fc# => X"9307c0fc",
		16#48fd# => X"635af700",
		16#48fe# => X"232a0100",
		16#48ff# => X"2328d100",
		16#4900# => X"13070000",
		16#4901# => X"6ff0dffb",
		16#4902# => X"8327c101",
		16#4903# => X"b7060800",
		16#4904# => X"93080000",
		16#4905# => X"b3e7d700",
		16#4906# => X"232ef100",
		16#4907# => X"9307d003",
		16#4908# => X"3387e740",
		16#4909# => X"13555740",
		16#490a# => X"93070300",
		16#490b# => X"1377f701",
		16#490c# => X"93060000",
		16#490d# => X"03a80700",
		16#490e# => X"93861600",
		16#490f# => X"93874700",
		16#4910# => X"b3e80801",
		16#4911# => X"e318d5fe",
		16#4912# => X"939e2600",
		16#4913# => X"631a0702",
		16#4914# => X"93073000",
		16#4915# => X"b387d740",
		16#4916# => X"63d8e700",
		16#4917# => X"93074000",
		16#4918# => X"b386d740",
		16#4919# => X"6f008006",
		16#491a# => X"3305d601",
		16#491b# => X"03250500",
		16#491c# => X"13071700",
		16#491d# => X"13064600",
		16#491e# => X"232ea6fe",
		16#491f# => X"6ff0dffd",
		16#4920# => X"93070102",
		16#4921# => X"b387d701",
		16#4922# => X"83a707ff",
		16#4923# => X"13080002",
		16#4924# => X"3308e840",
		16#4925# => X"b3970701",
		16#4926# => X"b3e8f800",
		16#4927# => X"93073000",
		16#4928# => X"130e0000",
		16#4929# => X"b387d740",
		16#492a# => X"6348fe04",
		16#492b# => X"13064000",
		16#492c# => X"b306d640",
		16#492d# => X"93972700",
		16#492e# => X"13060102",
		16#492f# => X"b307f600",
		16#4930# => X"0326c101",
		16#4931# => X"3357e600",
		16#4932# => X"23a8e7fe",
		16#4933# => X"13074000",
		16#4934# => X"93972600",
		16#4935# => X"b307f300",
		16#4936# => X"23a00700",
		16#4937# => X"93861600",
		16#4938# => X"e398e6fe",
		16#4939# => X"03270101",
		16#493a# => X"b3371001",
		16#493b# => X"b367f700",
		16#493c# => X"2328f100",
		16#493d# => X"6ff0dff0",
		16#493e# => X"330fd601",
		16#493f# => X"03250f00",
		16#4940# => X"032f4f00",
		16#4941# => X"130e1e00",
		16#4942# => X"3355e500",
		16#4943# => X"331f0f01",
		16#4944# => X"3365e501",
		16#4945# => X"2320a600",
		16#4946# => X"13064600",
		16#4947# => X"6ff0dff8",
		16#4948# => X"03264101",
		16#4949# => X"83278101",
		16#494a# => X"0328c101",
		16#494b# => X"b366f600",
		16#494c# => X"b3e60601",
		16#494d# => X"b3e6a600",
		16#494e# => X"63180700",
		16#494f# => X"b336d000",
		16#4950# => X"93070000",
		16#4951# => X"6ff05fe8",
		16#4952# => X"638a060c",
		16#4953# => X"9356c601",
		16#4954# => X"13184800",
		16#4955# => X"13964700",
		16#4956# => X"93d7c701",
		16#4957# => X"37074000",
		16#4958# => X"b3e6c600",
		16#4959# => X"b3e70701",
		16#495a# => X"b3e7e700",
		16#495b# => X"93f686ff",
		16#495c# => X"1307f07f",
		16#495d# => X"6ff05fe5",
		16#495e# => X"93070000",
		16#495f# => X"93060000",
		16#4960# => X"1307f07f",
		16#4961# => X"13968700",
		16#4962# => X"635e0600",
		16#4963# => X"13071700",
		16#4964# => X"1306f07f",
		16#4965# => X"6308c708",
		16#4966# => X"370680ff",
		16#4967# => X"1306f6ff",
		16#4968# => X"b3f7c700",
		16#4969# => X"1396d701",
		16#496a# => X"93d63600",
		16#496b# => X"b366d600",
		16#496c# => X"1306f07f",
		16#496d# => X"93d73700",
		16#496e# => X"631ec700",
		16#496f# => X"b3e6f600",
		16#4970# => X"93070000",
		16#4971# => X"63880600",
		16#4972# => X"b7070800",
		16#4973# => X"93060000",
		16#4974# => X"93050000",
		16#4975# => X"37061000",
		16#4976# => X"1306f6ff",
		16#4977# => X"b3f7c700",
		16#4978# => X"37061080",
		16#4979# => X"1377f77f",
		16#497a# => X"1306f6ff",
		16#497b# => X"13174701",
		16#497c# => X"b3f7c700",
		16#497d# => X"b3e7e700",
		16#497e# => X"37070080",
		16#497f# => X"1347f7ff",
		16#4980# => X"9395f501",
		16#4981# => X"b3f7e700",
		16#4982# => X"33e7b700",
		16#4983# => X"13850600",
		16#4984# => X"93050700",
		16#4985# => X"13010102",
		16#4986# => X"67800000",
		16#4987# => X"93070000",
		16#4988# => X"6ff01ff6",
		16#4989# => X"93070000",
		16#498a# => X"93060000",
		16#498b# => X"6ff09ff7",
		16#498c# => X"13060500",
		16#498d# => X"13050000",
		16#498e# => X"93f61500",
		16#498f# => X"63840600",
		16#4990# => X"3305c500",
		16#4991# => X"93d51500",
		16#4992# => X"13161600",
		16#4993# => X"e39605fe",
		16#4994# => X"67800000",
		16#4995# => X"63400506",
		16#4996# => X"63c60506",
		16#4997# => X"13860500",
		16#4998# => X"93050500",
		16#4999# => X"1305f0ff",
		16#499a# => X"630c0602",
		16#499b# => X"93061000",
		16#499c# => X"637ab600",
		16#499d# => X"6358c000",
		16#499e# => X"13161600",
		16#499f# => X"93961600",
		16#49a0# => X"e36ab6fe",
		16#49a1# => X"13050000",
		16#49a2# => X"63e6c500",
		16#49a3# => X"b385c540",
		16#49a4# => X"3365d500",
		16#49a5# => X"93d61600",
		16#49a6# => X"13561600",
		16#49a7# => X"e39606fe",
		16#49a8# => X"67800000",
		16#49a9# => X"93820000",
		16#49aa# => X"eff05ffb",
		16#49ab# => X"13850500",
		16#49ac# => X"67800200",
		16#49ad# => X"3305a040",
		16#49ae# => X"63d80500",
		16#49af# => X"b305b040",
		16#49b0# => X"6ff0dff9",
		16#49b1# => X"b305b040",
		16#49b2# => X"93820000",
		16#49b3# => X"eff01ff9",
		16#49b4# => X"3305a040",
		16#49b5# => X"67800200",
		16#49b6# => X"93820000",
		16#49b7# => X"63ca0500",
		16#49b8# => X"634c0500",
		16#49b9# => X"eff09ff7",
		16#49ba# => X"13850500",
		16#49bb# => X"67800200",
		16#49bc# => X"b305b040",
		16#49bd# => X"e35805fe",
		16#49be# => X"3305a040",
		16#49bf# => X"eff01ff6",
		16#49c0# => X"3305b040",
		16#49c1# => X"67800200",
		16#49c2# => X"b7070100",
		16#49c3# => X"637af502",
		16#49c4# => X"9307f00f",
		16#49c5# => X"b3b7a700",
		16#49c6# => X"93973700",
		16#49c7# => X"13070002",
		16#49c8# => X"3307f740",
		16#49c9# => X"b357f500",
		16#49ca# => X"37450110",
		16#49cb# => X"1305c56b",
		16#49cc# => X"b387a700",
		16#49cd# => X"03c50700",
		16#49ce# => X"3305a740",
		16#49cf# => X"67800000",
		16#49d0# => X"37070001",
		16#49d1# => X"93070001",
		16#49d2# => X"e36ae5fc",
		16#49d3# => X"93078001",
		16#49d4# => X"6ff0dffc",
		16#49d5# => X"130101ff",
		16#49d6# => X"13056000",
		16#49d7# => X"23261100",
		16#49d8# => X"ef000026",
		16#49d9# => X"13051000",
		16#49da# => X"efa0dfd1",
		16#49db# => X"03a5c181",
		16#49dc# => X"67800000",
		16#49dd# => X"130101ff",
		16#49de# => X"93050000",
		16#49df# => X"23248100",
		16#49e0# => X"23261100",
		16#49e1# => X"13040500",
		16#49e2# => X"ef00c02c",
		16#49e3# => X"03a58181",
		16#49e4# => X"8327c503",
		16#49e5# => X"63840700",
		16#49e6# => X"e7800700",
		16#49e7# => X"13050400",
		16#49e8# => X"efa05fce",
		16#49e9# => X"0327c52d",
		16#49ea# => X"63180704",
		16#49eb# => X"130101ff",
		16#49ec# => X"93050008",
		16#49ed# => X"23248100",
		16#49ee# => X"23261100",
		16#49ef# => X"13040500",
		16#49f0# => X"ef408fcf",
		16#49f1# => X"232ea42c",
		16#49f2# => X"9307f0ff",
		16#49f3# => X"630c0500",
		16#49f4# => X"93070508",
		16#49f5# => X"23200500",
		16#49f6# => X"13054500",
		16#49f7# => X"e31cf5fe",
		16#49f8# => X"93070000",
		16#49f9# => X"8320c100",
		16#49fa# => X"03248100",
		16#49fb# => X"13850700",
		16#49fc# => X"13010101",
		16#49fd# => X"67800000",
		16#49fe# => X"93070000",
		16#49ff# => X"13850700",
		16#4a00# => X"67800000",
		16#4a01# => X"130101ff",
		16#4a02# => X"23229100",
		16#4a03# => X"23261100",
		16#4a04# => X"23248100",
		16#4a05# => X"23202101",
		16#4a06# => X"1307f001",
		16#4a07# => X"93040500",
		16#4a08# => X"637ab700",
		16#4a09# => X"13076001",
		16#4a0a# => X"2320e500",
		16#4a0b# => X"1305f0ff",
		16#4a0c# => X"6f008002",
		16#4a0d# => X"8327c52d",
		16#4a0e# => X"13090600",
		16#4a0f# => X"13840500",
		16#4a10# => X"63880702",
		16#4a11# => X"93152400",
		16#4a12# => X"03a4c42d",
		16#4a13# => X"b305b400",
		16#4a14# => X"03a50500",
		16#4a15# => X"23a02501",
		16#4a16# => X"8320c100",
		16#4a17# => X"03248100",
		16#4a18# => X"83244100",
		16#4a19# => X"03290100",
		16#4a1a# => X"13010101",
		16#4a1b# => X"67800000",
		16#4a1c# => X"eff05ff3",
		16#4a1d# => X"e30805fc",
		16#4a1e# => X"6ff05ffb",
		16#4a1f# => X"9307f001",
		16#4a20# => X"63fab700",
		16#4a21# => X"93076001",
		16#4a22# => X"2320f500",
		16#4a23# => X"1305f0ff",
		16#4a24# => X"67800000",
		16#4a25# => X"8327c52d",
		16#4a26# => X"130101fe",
		16#4a27# => X"232c8100",
		16#4a28# => X"232e1100",
		16#4a29# => X"13860500",
		16#4a2a# => X"13040500",
		16#4a2b# => X"638a0700",
		16#4a2c# => X"13972500",
		16#4a2d# => X"b387e700",
		16#4a2e# => X"03a70700",
		16#4a2f# => X"63160702",
		16#4a30# => X"13050400",
		16#4a31# => X"2326c100",
		16#4a32# => X"ef008017",
		16#4a33# => X"93050500",
		16#4a34# => X"13050400",
		16#4a35# => X"03248101",
		16#4a36# => X"0326c100",
		16#4a37# => X"8320c101",
		16#4a38# => X"13010102",
		16#4a39# => X"6f00c010",
		16#4a3a# => X"93061000",
		16#4a3b# => X"13050000",
		16#4a3c# => X"630cd700",
		16#4a3d# => X"9306f0ff",
		16#4a3e# => X"6310d702",
		16#4a3f# => X"93076001",
		16#4a40# => X"2320f400",
		16#4a41# => X"13051000",
		16#4a42# => X"8320c101",
		16#4a43# => X"03248101",
		16#4a44# => X"13010102",
		16#4a45# => X"67800000",
		16#4a46# => X"13850500",
		16#4a47# => X"23a00700",
		16#4a48# => X"e7000700",
		16#4a49# => X"13050000",
		16#4a4a# => X"6ff01ffe",
		16#4a4b# => X"9307f001",
		16#4a4c# => X"63f6b700",
		16#4a4d# => X"1305f0ff",
		16#4a4e# => X"67800000",
		16#4a4f# => X"8327c52d",
		16#4a50# => X"130101ff",
		16#4a51# => X"23248100",
		16#4a52# => X"23229100",
		16#4a53# => X"23261100",
		16#4a54# => X"93040500",
		16#4a55# => X"13840500",
		16#4a56# => X"63840704",
		16#4a57# => X"83a7c42d",
		16#4a58# => X"13172400",
		16#4a59# => X"13051000",
		16#4a5a# => X"3387e700",
		16#4a5b# => X"83270700",
		16#4a5c# => X"638e0702",
		16#4a5d# => X"9306f0ff",
		16#4a5e# => X"13052000",
		16#4a5f# => X"6388d702",
		16#4a60# => X"93061000",
		16#4a61# => X"13053000",
		16#4a62# => X"6382d702",
		16#4a63# => X"13050400",
		16#4a64# => X"23200700",
		16#4a65# => X"e7800700",
		16#4a66# => X"13050000",
		16#4a67# => X"6f000001",
		16#4a68# => X"eff05fe0",
		16#4a69# => X"e30c05fa",
		16#4a6a# => X"1305f0ff",
		16#4a6b# => X"8320c100",
		16#4a6c# => X"03248100",
		16#4a6d# => X"83244100",
		16#4a6e# => X"13010101",
		16#4a6f# => X"67800000",
		16#4a70# => X"93050500",
		16#4a71# => X"03a5c181",
		16#4a72# => X"6ff05feb",
		16#4a73# => X"13860500",
		16#4a74# => X"93050500",
		16#4a75# => X"03a5c181",
		16#4a76# => X"6ff0dfe2",
		16#4a77# => X"03a5c181",
		16#4a78# => X"6ff05fdc",
		16#4a79# => X"93050500",
		16#4a7a# => X"03a5c181",
		16#4a7b# => X"6ff01ff4",
		16#4a7c# => X"130101ff",
		16#4a7d# => X"23248100",
		16#4a7e# => X"23229100",
		16#4a7f# => X"37840110",
		16#4a80# => X"93040500",
		16#4a81# => X"13850500",
		16#4a82# => X"93050600",
		16#4a83# => X"23261100",
		16#4a84# => X"232204aa",
		16#4a85# => X"efa0dfa4",
		16#4a86# => X"9307f0ff",
		16#4a87# => X"6318f500",
		16#4a88# => X"832744aa",
		16#4a89# => X"63840700",
		16#4a8a# => X"23a0f400",
		16#4a8b# => X"8320c100",
		16#4a8c# => X"03248100",
		16#4a8d# => X"83244100",
		16#4a8e# => X"13010101",
		16#4a8f# => X"67800000",
		16#4a90# => X"6fa09fa1",
		16#4a91# => X"13860500",
		16#4a92# => X"93050500",
		16#4a93# => X"03a5c181",
		16#4a94# => X"6ff01ffa",
		16#4a95# => X"130101fd",
		16#4a96# => X"232e3101",
		16#4a97# => X"83a98181",
		16#4a98# => X"232c4101",
		16#4a99# => X"232a5101",
		16#4a9a# => X"23286101",
		16#4a9b# => X"23261102",
		16#4a9c# => X"23248102",
		16#4a9d# => X"23229102",
		16#4a9e# => X"23202103",
		16#4a9f# => X"23267101",
		16#4aa0# => X"930a0500",
		16#4aa1# => X"138a0500",
		16#4aa2# => X"130b1000",
		16#4aa3# => X"83a48914",
		16#4aa4# => X"638c0400",
		16#4aa5# => X"03a44400",
		16#4aa6# => X"1309f4ff",
		16#4aa7# => X"13142400",
		16#4aa8# => X"33848400",
		16#4aa9# => X"63580902",
		16#4aaa# => X"8320c102",
		16#4aab# => X"03248102",
		16#4aac# => X"83244102",
		16#4aad# => X"03290102",
		16#4aae# => X"8329c101",
		16#4aaf# => X"032a8101",
		16#4ab0# => X"832a4101",
		16#4ab1# => X"032b0101",
		16#4ab2# => X"832bc100",
		16#4ab3# => X"13010103",
		16#4ab4# => X"67800000",
		16#4ab5# => X"630c0a00",
		16#4ab6# => X"83274410",
		16#4ab7# => X"63884701",
		16#4ab8# => X"1309f9ff",
		16#4ab9# => X"1304c4ff",
		16#4aba# => X"6ff0dffb",
		16#4abb# => X"03a74400",
		16#4abc# => X"83274400",
		16#4abd# => X"1307f7ff",
		16#4abe# => X"631c2703",
		16#4abf# => X"23a22401",
		16#4ac0# => X"e38007fe",
		16#4ac1# => X"83a68418",
		16#4ac2# => X"33172b01",
		16#4ac3# => X"83ab4400",
		16#4ac4# => X"b376d700",
		16#4ac5# => X"63920602",
		16#4ac6# => X"e7800700",
		16#4ac7# => X"03a74400",
		16#4ac8# => X"83a78914",
		16#4ac9# => X"e31477f7",
		16#4aca# => X"e38cf4fa",
		16#4acb# => X"6ff01ff6",
		16#4acc# => X"23220400",
		16#4acd# => X"6ff0dffc",
		16#4ace# => X"83a6c418",
		16#4acf# => X"83254408",
		16#4ad0# => X"3377d700",
		16#4ad1# => X"63180700",
		16#4ad2# => X"13850a00",
		16#4ad3# => X"e7800700",
		16#4ad4# => X"6ff0dffc",
		16#4ad5# => X"13850500",
		16#4ad6# => X"e7800700",
		16#4ad7# => X"6ff01ffc",
		16#4ad8# => X"130101f6",
		16#4ad9# => X"232e1108",
		16#4ada# => X"232c8108",
		16#4adb# => X"2326b107",
		16#4adc# => X"1304010a",
		16#4add# => X"232a9108",
		16#4ade# => X"23282109",
		16#4adf# => X"23263109",
		16#4ae0# => X"23244109",
		16#4ae1# => X"23225109",
		16#4ae2# => X"23206109",
		16#4ae3# => X"232e7107",
		16#4ae4# => X"232c8107",
		16#4ae5# => X"232a9107",
		16#4ae6# => X"2328a107",
		16#4ae7# => X"b7370110",
		16#4ae8# => X"83a30734",
		16#4ae9# => X"130101fc",
		16#4aea# => X"13870734",
		16#4aeb# => X"13060100",
		16#4aec# => X"b7460110",
		16#4aed# => X"130101fc",
		16#4aee# => X"93874689",
		16#4aef# => X"832f8700",
		16#4af0# => X"032fc700",
		16#4af1# => X"832e0701",
		16#4af2# => X"032e4701",
		16#4af3# => X"03238701",
		16#4af4# => X"83224700",
		16#4af5# => X"8358c701",
		16#4af6# => X"0348e701",
		16#4af7# => X"83a54689",
		16#4af8# => X"13072000",
		16#4af9# => X"93060100",
		16#4afa# => X"23a4e600",
		16#4afb# => X"23a87600",
		16#4afc# => X"13078002",
		16#4afd# => X"b7830110",
		16#4afe# => X"b78d0110",
		16#4aff# => X"23a2c39c",
		16#4b00# => X"23a0c600",
		16#4b01# => X"23a6e600",
		16#4b02# => X"23a20600",
		16#4b03# => X"23a8dd9c",
		16#4b04# => X"03a54700",
		16#4b05# => X"23aa5600",
		16#4b06# => X"03d7c701",
		16#4b07# => X"03a64701",
		16#4b08# => X"23acf601",
		16#4b09# => X"23aee601",
		16#4b0a# => X"23a0d603",
		16#4b0b# => X"23a2c603",
		16#4b0c# => X"23a46602",
		16#4b0d# => X"23961603",
		16#4b0e# => X"23870603",
		16#4b0f# => X"83a88700",
		16#4b10# => X"03a8c700",
		16#4b11# => X"83a68701",
		16#4b12# => X"2320b4f8",
		16#4b13# => X"83a50701",
		16#4b14# => X"83c7e701",
		16#4b15# => X"231ee4f8",
		16#4b16# => X"37570110",
		16#4b17# => X"1307072b",
		16#4b18# => X"2322a4f8",
		16#4b19# => X"230ff4f8",
		16#4b1a# => X"1305a000",
		16#4b1b# => X"9307a000",
		16#4b1c# => X"232ef764",
		16#4b1d# => X"232414f9",
		16#4b1e# => X"232604f9",
		16#4b1f# => X"2328b4f8",
		16#4b20# => X"232ac4f8",
		16#4b21# => X"232cd4f8",
		16#4b22# => X"efe0de88",
		16#4b23# => X"b7350110",
		16#4b24# => X"37350110",
		16#4b25# => X"93850536",
		16#4b26# => X"13050537",
		16#4b27# => X"efe05e82",
		16#4b28# => X"b7570110",
		16#4b29# => X"83a7c724",
		16#4b2a# => X"63820766",
		16#4b2b# => X"37350110",
		16#4b2c# => X"13054539",
		16#4b2d# => X"efe09e9d",
		16#4b2e# => X"b7350110",
		16#4b2f# => X"37350110",
		16#4b30# => X"13061000",
		16#4b31# => X"9385053f",
		16#4b32# => X"1305853f",
		16#4b33# => X"efe04eff",
		16#4b34# => X"1305a000",
		16#4b35# => X"efe01e84",
		16#4b36# => X"374a0110",
		16#4b37# => X"83274a8b",
		16#4b38# => X"378b0110",
		16#4b39# => X"130a4a8b",
		16#4b3a# => X"2326f4f6",
		16#4b3b# => X"b7470110",
		16#4b3c# => X"83ac478d",
		16#4b3d# => X"b7870110",
		16#4b3e# => X"23aa079c",
		16#4b3f# => X"9307a000",
		16#4b40# => X"2324f4f6",
		16#4b41# => X"378c0110",
		16#4b42# => X"032984f6",
		16#4b43# => X"b7370110",
		16#4b44# => X"1385c740",
		16#4b45# => X"93050900",
		16#4b46# => X"efe08efa",
		16#4b47# => X"13858187",
		16#4b48# => X"93840700",
		16#4b49# => X"efe0deb0",
		16#4b4a# => X"83a78187",
		16#4b4b# => X"130d1900",
		16#4b4c# => X"930b1000",
		16#4b4d# => X"23aaf188",
		16#4b4e# => X"930a2000",
		16#4b4f# => X"efe0cef2",
		16#4b50# => X"efe08eef",
		16#4b51# => X"8347ea01",
		16#4b52# => X"03264a01",
		16#4b53# => X"032e4a00",
		16#4b54# => X"03238a00",
		16#4b55# => X"8328ca00",
		16#4b56# => X"03280a01",
		16#4b57# => X"83268a01",
		16#4b58# => X"0357ca01",
		16#4b59# => X"832ec4f6",
		16#4b5a# => X"230ff4fa",
		16#4b5b# => X"930504fa",
		16#4b5c# => X"93071000",
		16#4b5d# => X"130504f8",
		16#4b5e# => X"232ac4fa",
		16#4b5f# => X"232ef4f6",
		16#4b60# => X"232a54f7",
		16#4b61# => X"2320d4fb",
		16#4b62# => X"2322c4fb",
		16#4b63# => X"232464fa",
		16#4b64# => X"232614fb",
		16#4b65# => X"232804fb",
		16#4b66# => X"232cd4fa",
		16#4b67# => X"231ee4fa",
		16#4b68# => X"efe00eb8",
		16#4b69# => X"032644f7",
		16#4b6a# => X"13351500",
		16#4b6b# => X"b7870110",
		16#4b6c# => X"23a0a7aa",
		16#4b6d# => X"63ccca02",
		16#4b6e# => X"13050600",
		16#4b6f# => X"93172500",
		16#4b70# => X"b387a700",
		16#4b71# => X"9387d7ff",
		16#4b72# => X"130684f7",
		16#4b73# => X"93053000",
		16#4b74# => X"232cf4f6",
		16#4b75# => X"efe04ea7",
		16#4b76# => X"032544f7",
		16#4b77# => X"13051500",
		16#4b78# => X"232aa4f6",
		16#4b79# => X"e3dcaafc",
		16#4b7a# => X"13060500",
		16#4b7b# => X"832684f7",
		16#4b7c# => X"b7570110",
		16#4b7d# => X"9385072b",
		16#4b7e# => X"b7870110",
		16#4b7f# => X"1385879d",
		16#4b80# => X"efe08ea5",
		16#4b81# => X"03a50d9d",
		16#4b82# => X"efe00ecd",
		16#4b83# => X"0347db9c",
		16#4b84# => X"93070004",
		16#4b85# => X"63fce74a",
		16#4b86# => X"b7470110",
		16#4b87# => X"13091004",
		16#4b88# => X"93093000",
		16#4b89# => X"9384478d",
		16#4b8a# => X"6f004001",
		16#4b8b# => X"8347db9c",
		16#4b8c# => X"13091900",
		16#4b8d# => X"1379f90f",
		16#4b8e# => X"63e02709",
		16#4b8f# => X"93053004",
		16#4b90# => X"13050900",
		16#4b91# => X"efe08eab",
		16#4b92# => X"8327c4f7",
		16#4b93# => X"e310f5fe",
		16#4b94# => X"9305c4f7",
		16#4b95# => X"13050000",
		16#4b96# => X"efe08eb3",
		16#4b97# => X"83c7e401",
		16#4b98# => X"83a84400",
		16#4b99# => X"03a88400",
		16#4b9a# => X"03a5c400",
		16#4b9b# => X"83a50401",
		16#4b9c# => X"03a64401",
		16#4b9d# => X"83a68401",
		16#4b9e# => X"03d7c401",
		16#4b9f# => X"230ff4fa",
		16#4ba0# => X"8347db9c",
		16#4ba1# => X"13091900",
		16#4ba2# => X"232094fb",
		16#4ba3# => X"232214fb",
		16#4ba4# => X"232404fb",
		16#4ba5# => X"2326a4fa",
		16#4ba6# => X"2328b4fa",
		16#4ba7# => X"232ac4fa",
		16#4ba8# => X"232cd4fa",
		16#4ba9# => X"231ee4fa",
		16#4baa# => X"23247c9d",
		16#4bab# => X"1379f90f",
		16#4bac# => X"93890b00",
		16#4bad# => X"e3f427f9",
		16#4bae# => X"832544f7",
		16#4baf# => X"13850900",
		16#4bb0# => X"938b1b00",
		16#4bb1# => X"eff0cff6",
		16#4bb2# => X"032984f7",
		16#4bb3# => X"93090500",
		16#4bb4# => X"93050900",
		16#4bb5# => X"eff00ff8",
		16#4bb6# => X"93040500",
		16#4bb7# => X"130544f7",
		16#4bb8# => X"232a94f6",
		16#4bb9# => X"efe08eb9",
		16#4bba# => X"e39aabe5",
		16#4bbb# => X"13858187",
		16#4bbc# => X"938a0700",
		16#4bbd# => X"efe0de93",
		16#4bbe# => X"83a58187",
		16#4bbf# => X"83a74189",
		16#4bc0# => X"37870110",
		16#4bc1# => X"2320b79c",
		16#4bc2# => X"b385f540",
		16#4bc3# => X"23a8b188",
		16#4bc4# => X"6352b03c",
		16#4bc5# => X"93071000",
		16#4bc6# => X"37870110",
		16#4bc7# => X"232af79c",
		16#4bc8# => X"37350110",
		16#4bc9# => X"1305c546",
		16#4bca# => X"efe04ef6",
		16#4bcb# => X"1305a000",
		16#4bcc# => X"efe04ede",
		16#4bcd# => X"83258c9c",
		16#4bce# => X"37350110",
		16#4bcf# => X"1305454a",
		16#4bd0# => X"373a0110",
		16#4bd1# => X"efe0ced7",
		16#4bd2# => X"93055000",
		16#4bd3# => X"13050a4c",
		16#4bd4# => X"efe00ed7",
		16#4bd5# => X"b7870110",
		16#4bd6# => X"83a507aa",
		16#4bd7# => X"37350110",
		16#4bd8# => X"1305c54d",
		16#4bd9# => X"efe0ced5",
		16#4bda# => X"93051000",
		16#4bdb# => X"13050a4c",
		16#4bdc# => X"efe00ed5",
		16#4bdd# => X"b7870110",
		16#4bde# => X"83c5c79c",
		16#4bdf# => X"37350110",
		16#4be0# => X"1305854f",
		16#4be1# => X"efe0ced3",
		16#4be2# => X"b73a0110",
		16#4be3# => X"93051004",
		16#4be4# => X"13854a51",
		16#4be5# => X"efe0ced2",
		16#4be6# => X"8345db9c",
		16#4be7# => X"37350110",
		16#4be8# => X"13050553",
		16#4be9# => X"efe0ced1",
		16#4bea# => X"93052004",
		16#4beb# => X"13854a51",
		16#4bec# => X"efe00ed1",
		16#4bed# => X"b7870110",
		16#4bee# => X"9387879d",
		16#4bef# => X"83a50702",
		16#4bf0# => X"37350110",
		16#4bf1# => X"1305c554",
		16#4bf2# => X"efe08ecf",
		16#4bf3# => X"93057000",
		16#4bf4# => X"13050a4c",
		16#4bf5# => X"efe0cece",
		16#4bf6# => X"b7570110",
		16#4bf7# => X"9387072b",
		16#4bf8# => X"83a5c765",
		16#4bf9# => X"37350110",
		16#4bfa# => X"13058556",
		16#4bfb# => X"efe04ecd",
		16#4bfc# => X"37350110",
		16#4bfd# => X"13054558",
		16#4bfe# => X"efe04ee9",
		16#4bff# => X"37350110",
		16#4c00# => X"1305055b",
		16#4c01# => X"efe08ee8",
		16#4c02# => X"03a70d9d",
		16#4c03# => X"b7370110",
		16#4c04# => X"1385c75b",
		16#4c05# => X"83250700",
		16#4c06# => X"2326f4f6",
		16#4c07# => X"373d0110",
		16#4c08# => X"efe00eca",
		16#4c09# => X"37350110",
		16#4c0a# => X"1305855d",
		16#4c0b# => X"efe00ee6",
		16#4c0c# => X"03a70d9d",
		16#4c0d# => X"b7370110",
		16#4c0e# => X"13858760",
		16#4c0f# => X"83254700",
		16#4c10# => X"b73c0110",
		16#4c11# => X"373c0110",
		16#4c12# => X"efe08ec7",
		16#4c13# => X"93050000",
		16#4c14# => X"13050a4c",
		16#4c15# => X"efe0cec6",
		16#4c16# => X"03a70d9d",
		16#4c17# => X"13054d62",
		16#4c18# => X"b73b0110",
		16#4c19# => X"83258700",
		16#4c1a# => X"33892941",
		16#4c1b# => X"efe04ec5",
		16#4c1c# => X"93052000",
		16#4c1d# => X"13050a4c",
		16#4c1e# => X"efe08ec4",
		16#4c1f# => X"03a70d9d",
		16#4c20# => X"13850c64",
		16#4c21# => X"8325c700",
		16#4c22# => X"efe08ec3",
		16#4c23# => X"93051001",
		16#4c24# => X"13050a4c",
		16#4c25# => X"efe0cec2",
		16#4c26# => X"83a50d9d",
		16#4c27# => X"1305cc65",
		16#4c28# => X"b78d0110",
		16#4c29# => X"93850501",
		16#4c2a# => X"efe08ec1",
		16#4c2b# => X"13858b67",
		16#4c2c# => X"efe0cedd",
		16#4c2d# => X"37350110",
		16#4c2e# => X"1305c56a",
		16#4c2f# => X"efe00edd",
		16#4c30# => X"03a74d9c",
		16#4c31# => X"8327c4f6",
		16#4c32# => X"83250700",
		16#4c33# => X"1385c75b",
		16#4c34# => X"efe00ebf",
		16#4c35# => X"37350110",
		16#4c36# => X"1305c56b",
		16#4c37# => X"efe00edb",
		16#4c38# => X"83a74d9c",
		16#4c39# => X"37370110",
		16#4c3a# => X"13058760",
		16#4c3b# => X"83a54700",
		16#4c3c# => X"efe00ebd",
		16#4c3d# => X"93050000",
		16#4c3e# => X"13050a4c",
		16#4c3f# => X"efe04ebc",
		16#4c40# => X"83a74d9c",
		16#4c41# => X"13054d62",
		16#4c42# => X"83a58700",
		16#4c43# => X"efe04ebb",
		16#4c44# => X"93051000",
		16#4c45# => X"13050a4c",
		16#4c46# => X"efe08eba",
		16#4c47# => X"83a74d9c",
		16#4c48# => X"13850c64",
		16#4c49# => X"83a5c700",
		16#4c4a# => X"efe08eb9",
		16#4c4b# => X"93052001",
		16#4c4c# => X"13050a4c",
		16#4c4d# => X"efe0ceb8",
		16#4c4e# => X"83a54d9c",
		16#4c4f# => X"1305cc65",
		16#4c50# => X"93850501",
		16#4c51# => X"efe0ceb7",
		16#4c52# => X"13858b67",
		16#4c53# => X"efe00ed4",
		16#4c54# => X"832544f7",
		16#4c55# => X"37350110",
		16#4c56# => X"1305c56f",
		16#4c57# => X"efe04eb6",
		16#4c58# => X"93055000",
		16#4c59# => X"13050a4c",
		16#4c5a# => X"efe08eb5",
		16#4c5b# => X"93173900",
		16#4c5c# => X"33892741",
		16#4c5d# => X"37350110",
		16#4c5e# => X"b3059940",
		16#4c5f# => X"13058571",
		16#4c60# => X"efe00eb4",
		16#4c61# => X"9305d000",
		16#4c62# => X"13050a4c",
		16#4c63# => X"efe04eb3",
		16#4c64# => X"832584f7",
		16#4c65# => X"37350110",
		16#4c66# => X"13054573",
		16#4c67# => X"efe04eb2",
		16#4c68# => X"93057000",
		16#4c69# => X"13050a4c",
		16#4c6a# => X"efe08eb1",
		16#4c6b# => X"8325c4f7",
		16#4c6c# => X"37350110",
		16#4c6d# => X"13050575",
		16#4c6e# => X"efe08eb0",
		16#4c6f# => X"93051000",
		16#4c70# => X"13050a4c",
		16#4c71# => X"efe0ceaf",
		16#4c72# => X"37350110",
		16#4c73# => X"930504f8",
		16#4c74# => X"1305c576",
		16#4c75# => X"efe0ceae",
		16#4c76# => X"37350110",
		16#4c77# => X"13058578",
		16#4c78# => X"efe0ceca",
		16#4c79# => X"37350110",
		16#4c7a# => X"930504fa",
		16#4c7b# => X"1305c57b",
		16#4c7c# => X"efe00ead",
		16#4c7d# => X"37350110",
		16#4c7e# => X"1305857d",
		16#4c7f# => X"efe00ec9",
		16#4c80# => X"1305a000",
		16#4c81# => X"efe00eb1",
		16#4c82# => X"83a40189",
		16#4c83# => X"b7450f00",
		16#4c84# => X"93850524",
		16#4c85# => X"13850400",
		16#4c86# => X"eff08fc1",
		16#4c87# => X"832984f6",
		16#4c88# => X"93850900",
		16#4c89# => X"eff00fc3",
		16#4c8a# => X"13090500",
		16#4c8b# => X"93850400",
		16#4c8c# => X"23a4a188",
		16#4c8d# => X"13850900",
		16#4c8e# => X"eff0cfc1",
		16#4c8f# => X"23a6a188",
		16#4c90# => X"93050900",
		16#4c91# => X"13850400",
		16#4c92# => X"eff08fbe",
		16#4c93# => X"93850900",
		16#4c94# => X"eff04fc0",
		16#4c95# => X"13060500",
		16#4c96# => X"37450110",
		16#4c97# => X"93850400",
		16#4c98# => X"1305c580",
		16#4c99# => X"efe0cea5",
		16#4c9a# => X"83a58188",
		16#4c9b# => X"37450110",
		16#4c9c# => X"1305c582",
		16#4c9d# => X"efe0cea4",
		16#4c9e# => X"83a5c188",
		16#4c9f# => X"37450110",
		16#4ca0# => X"13050586",
		16#4ca1# => X"efe0cea3",
		16#4ca2# => X"130104f6",
		16#4ca3# => X"8320c109",
		16#4ca4# => X"13050000",
		16#4ca5# => X"03248109",
		16#4ca6# => X"83244109",
		16#4ca7# => X"03290109",
		16#4ca8# => X"8329c108",
		16#4ca9# => X"032a8108",
		16#4caa# => X"832a4108",
		16#4cab# => X"032b0108",
		16#4cac# => X"832bc107",
		16#4cad# => X"032c8107",
		16#4cae# => X"832c4107",
		16#4caf# => X"032d0107",
		16#4cb0# => X"832dc106",
		16#4cb1# => X"1301010a",
		16#4cb2# => X"67800000",
		16#4cb3# => X"93093000",
		16#4cb4# => X"6ff09fbe",
		16#4cb5# => X"37350110",
		16#4cb6# => X"13050543",
		16#4cb7# => X"efe04e9e",
		16#4cb8# => X"032784f6",
		16#4cb9# => X"1305a000",
		16#4cba# => X"93172700",
		16#4cbb# => X"b387e700",
		16#4cbc# => X"93971700",
		16#4cbd# => X"2324f4f6",
		16#4cbe# => X"efe0cea1",
		16#4cbf# => X"b7870110",
		16#4cc0# => X"83a7479d",
		16#4cc1# => X"e38207a0",
		16#4cc2# => X"6ff09fc1",
		16#4cc3# => X"37350110",
		16#4cc4# => X"1305053c",
		16#4cc5# => X"efe08eb7",
		16#4cc6# => X"6ff01f9a",
		16#4cc7# => X"37450110",
		16#4cc8# => X"130101ff",
		16#4cc9# => X"13058596",
		16#4cca# => X"23261100",
		16#4ccb# => X"efe00eb6",
		16#4ccc# => X"8320c100",
		16#4ccd# => X"1305f0ff",
		16#4cce# => X"13010101",
		16#4ccf# => X"67800000",
		16#4cd0# => X"44485259",
		16#4cd1# => X"53544f4e",
		16#4cd2# => X"45205052",
		16#4cd3# => X"4f475241",
		16#4cd4# => X"4d2c2053",
		16#4cd5# => X"4f4d4520",
		16#4cd6# => X"53545249",
		16#4cd7# => X"4e470000",
		16#4cd8# => X"432c2056",
		16#4cd9# => X"65727369",
		16#4cda# => X"6f6e2032",
		16#4cdb# => X"2e320000",
		16#4cdc# => X"44687279",
		16#4cdd# => X"73746f6e",
		16#4cde# => X"65204265",
		16#4cdf# => X"6e63686d",
		16#4ce0# => X"61726b2c",
		16#4ce1# => X"20566572",
		16#4ce2# => X"73696f6e",
		16#4ce3# => X"2025730a",
		16#4ce4# => X"00000000",
		16#4ce5# => X"50726f67",
		16#4ce6# => X"72616d20",
		16#4ce7# => X"636f6d70",
		16#4ce8# => X"696c6564",
		16#4ce9# => X"20776974",
		16#4cea# => X"68202772",
		16#4ceb# => X"65676973",
		16#4cec# => X"74657227",
		16#4ced# => X"20617474",
		16#4cee# => X"72696275",
		16#4cef# => X"74650000",
		16#4cf0# => X"50726f67",
		16#4cf1# => X"72616d20",
		16#4cf2# => X"636f6d70",
		16#4cf3# => X"696c6564",
		16#4cf4# => X"20776974",
		16#4cf5# => X"686f7574",
		16#4cf6# => X"20277265",
		16#4cf7# => X"67697374",
		16#4cf8# => X"65722720",
		16#4cf9# => X"61747472",
		16#4cfa# => X"69627574",
		16#4cfb# => X"65000000",
		16#4cfc# => X"74696d65",
		16#4cfd# => X"73282900",
		16#4cfe# => X"5573696e",
		16#4cff# => X"67202573",
		16#4d00# => X"2c20485a",
		16#4d01# => X"3d25640a",
		16#4d02# => X"00000000",
		16#4d03# => X"54727969",
		16#4d04# => X"6e672025",
		16#4d05# => X"64207275",
		16#4d06# => X"6e732074",
		16#4d07# => X"68726f75",
		16#4d08# => X"67682044",
		16#4d09# => X"68727973",
		16#4d0a# => X"746f6e65",
		16#4d0b# => X"3a0a0000",
		16#4d0c# => X"4d656173",
		16#4d0d# => X"75726564",
		16#4d0e# => X"2074696d",
		16#4d0f# => X"6520746f",
		16#4d10# => X"6f20736d",
		16#4d11# => X"616c6c20",
		16#4d12# => X"746f206f",
		16#4d13# => X"62746169",
		16#4d14# => X"6e206d65",
		16#4d15# => X"616e696e",
		16#4d16# => X"6766756c",
		16#4d17# => X"20726573",
		16#4d18# => X"756c7473",
		16#4d19# => X"3a202564",
		16#4d1a# => X"0a000000",
		16#4d1b# => X"46696e61",
		16#4d1c# => X"6c207661",
		16#4d1d# => X"6c756573",
		16#4d1e# => X"206f6620",
		16#4d1f# => X"74686520",
		16#4d20# => X"76617269",
		16#4d21# => X"61626c65",
		16#4d22# => X"73207573",
		16#4d23# => X"65642069",
		16#4d24# => X"6e207468",
		16#4d25# => X"65206265",
		16#4d26# => X"6e63686d",
		16#4d27# => X"61726b3a",
		16#4d28# => X"00000000",
		16#4d29# => X"496e745f",
		16#4d2a# => X"476c6f62",
		16#4d2b# => X"3a202020",
		16#4d2c# => X"20202020",
		16#4d2d# => X"20202020",
		16#4d2e# => X"2025640a",
		16#4d2f# => X"00000000",
		16#4d30# => X"20202020",
		16#4d31# => X"20202020",
		16#4d32# => X"73686f75",
		16#4d33# => X"6c642062",
		16#4d34# => X"653a2020",
		16#4d35# => X"2025640a",
		16#4d36# => X"00000000",
		16#4d37# => X"426f6f6c",
		16#4d38# => X"5f476c6f",
		16#4d39# => X"623a2020",
		16#4d3a# => X"20202020",
		16#4d3b# => X"20202020",
		16#4d3c# => X"2025640a",
		16#4d3d# => X"00000000",
		16#4d3e# => X"43685f31",
		16#4d3f# => X"5f476c6f",
		16#4d40# => X"623a2020",
		16#4d41# => X"20202020",
		16#4d42# => X"20202020",
		16#4d43# => X"2025630a",
		16#4d44# => X"00000000",
		16#4d45# => X"20202020",
		16#4d46# => X"20202020",
		16#4d47# => X"73686f75",
		16#4d48# => X"6c642062",
		16#4d49# => X"653a2020",
		16#4d4a# => X"2025630a",
		16#4d4b# => X"00000000",
		16#4d4c# => X"43685f32",
		16#4d4d# => X"5f476c6f",
		16#4d4e# => X"623a2020",
		16#4d4f# => X"20202020",
		16#4d50# => X"20202020",
		16#4d51# => X"2025630a",
		16#4d52# => X"00000000",
		16#4d53# => X"4172725f",
		16#4d54# => X"315f476c",
		16#4d55# => X"6f625b38",
		16#4d56# => X"5d3a2020",
		16#4d57# => X"20202020",
		16#4d58# => X"2025640a",
		16#4d59# => X"00000000",
		16#4d5a# => X"4172725f",
		16#4d5b# => X"325f476c",
		16#4d5c# => X"6f625b38",
		16#4d5d# => X"5d5b375d",
		16#4d5e# => X"3a202020",
		16#4d5f# => X"2025640a",
		16#4d60# => X"00000000",
		16#4d61# => X"20202020",
		16#4d62# => X"20202020",
		16#4d63# => X"73686f75",
		16#4d64# => X"6c642062",
		16#4d65# => X"653a2020",
		16#4d66# => X"204e756d",
		16#4d67# => X"6265725f",
		16#4d68# => X"4f665f52",
		16#4d69# => X"756e7320",
		16#4d6a# => X"2b203130",
		16#4d6b# => X"00000000",
		16#4d6c# => X"5074725f",
		16#4d6d# => X"476c6f62",
		16#4d6e# => X"2d3e0000",
		16#4d6f# => X"20205074",
		16#4d70# => X"725f436f",
		16#4d71# => X"6d703a20",
		16#4d72# => X"20202020",
		16#4d73# => X"20202020",
		16#4d74# => X"2025640a",
		16#4d75# => X"00000000",
		16#4d76# => X"20202020",
		16#4d77# => X"20202020",
		16#4d78# => X"73686f75",
		16#4d79# => X"6c642062",
		16#4d7a# => X"653a2020",
		16#4d7b# => X"2028696d",
		16#4d7c# => X"706c656d",
		16#4d7d# => X"656e7461",
		16#4d7e# => X"74696f6e",
		16#4d7f# => X"2d646570",
		16#4d80# => X"656e6465",
		16#4d81# => X"6e742900",
		16#4d82# => X"20204469",
		16#4d83# => X"7363723a",
		16#4d84# => X"20202020",
		16#4d85# => X"20202020",
		16#4d86# => X"20202020",
		16#4d87# => X"2025640a",
		16#4d88# => X"00000000",
		16#4d89# => X"2020456e",
		16#4d8a# => X"756d5f43",
		16#4d8b# => X"6f6d703a",
		16#4d8c# => X"20202020",
		16#4d8d# => X"20202020",
		16#4d8e# => X"2025640a",
		16#4d8f# => X"00000000",
		16#4d90# => X"2020496e",
		16#4d91# => X"745f436f",
		16#4d92# => X"6d703a20",
		16#4d93# => X"20202020",
		16#4d94# => X"20202020",
		16#4d95# => X"2025640a",
		16#4d96# => X"00000000",
		16#4d97# => X"20205374",
		16#4d98# => X"725f436f",
		16#4d99# => X"6d703a20",
		16#4d9a# => X"20202020",
		16#4d9b# => X"20202020",
		16#4d9c# => X"2025730a",
		16#4d9d# => X"00000000",
		16#4d9e# => X"20202020",
		16#4d9f# => X"20202020",
		16#4da0# => X"73686f75",
		16#4da1# => X"6c642062",
		16#4da2# => X"653a2020",
		16#4da3# => X"20444852",
		16#4da4# => X"5953544f",
		16#4da5# => X"4e452050",
		16#4da6# => X"524f4752",
		16#4da7# => X"414d2c20",
		16#4da8# => X"534f4d45",
		16#4da9# => X"20535452",
		16#4daa# => X"494e4700",
		16#4dab# => X"4e657874",
		16#4dac# => X"5f507472",
		16#4dad# => X"5f476c6f",
		16#4dae# => X"622d3e00",
		16#4daf# => X"20202020",
		16#4db0# => X"20202020",
		16#4db1# => X"73686f75",
		16#4db2# => X"6c642062",
		16#4db3# => X"653a2020",
		16#4db4# => X"2028696d",
		16#4db5# => X"706c656d",
		16#4db6# => X"656e7461",
		16#4db7# => X"74696f6e",
		16#4db8# => X"2d646570",
		16#4db9# => X"656e6465",
		16#4dba# => X"6e74292c",
		16#4dbb# => X"2073616d",
		16#4dbc# => X"65206173",
		16#4dbd# => X"2061626f",
		16#4dbe# => X"76650000",
		16#4dbf# => X"496e745f",
		16#4dc0# => X"315f4c6f",
		16#4dc1# => X"633a2020",
		16#4dc2# => X"20202020",
		16#4dc3# => X"20202020",
		16#4dc4# => X"2025640a",
		16#4dc5# => X"00000000",
		16#4dc6# => X"496e745f",
		16#4dc7# => X"325f4c6f",
		16#4dc8# => X"633a2020",
		16#4dc9# => X"20202020",
		16#4dca# => X"20202020",
		16#4dcb# => X"2025640a",
		16#4dcc# => X"00000000",
		16#4dcd# => X"496e745f",
		16#4dce# => X"335f4c6f",
		16#4dcf# => X"633a2020",
		16#4dd0# => X"20202020",
		16#4dd1# => X"20202020",
		16#4dd2# => X"2025640a",
		16#4dd3# => X"00000000",
		16#4dd4# => X"456e756d",
		16#4dd5# => X"5f4c6f63",
		16#4dd6# => X"3a202020",
		16#4dd7# => X"20202020",
		16#4dd8# => X"20202020",
		16#4dd9# => X"2025640a",
		16#4dda# => X"00000000",
		16#4ddb# => X"5374725f",
		16#4ddc# => X"315f4c6f",
		16#4ddd# => X"633a2020",
		16#4dde# => X"20202020",
		16#4ddf# => X"20202020",
		16#4de0# => X"2025730a",
		16#4de1# => X"00000000",
		16#4de2# => X"20202020",
		16#4de3# => X"20202020",
		16#4de4# => X"73686f75",
		16#4de5# => X"6c642062",
		16#4de6# => X"653a2020",
		16#4de7# => X"20444852",
		16#4de8# => X"5953544f",
		16#4de9# => X"4e452050",
		16#4dea# => X"524f4752",
		16#4deb# => X"414d2c20",
		16#4dec# => X"31275354",
		16#4ded# => X"20535452",
		16#4dee# => X"494e4700",
		16#4def# => X"5374725f",
		16#4df0# => X"325f4c6f",
		16#4df1# => X"633a2020",
		16#4df2# => X"20202020",
		16#4df3# => X"20202020",
		16#4df4# => X"2025730a",
		16#4df5# => X"00000000",
		16#4df6# => X"20202020",
		16#4df7# => X"20202020",
		16#4df8# => X"73686f75",
		16#4df9# => X"6c642062",
		16#4dfa# => X"653a2020",
		16#4dfb# => X"20444852",
		16#4dfc# => X"5953544f",
		16#4dfd# => X"4e452050",
		16#4dfe# => X"524f4752",
		16#4dff# => X"414d2c20",
		16#4e00# => X"32274e44",
		16#4e01# => X"20535452",
		16#4e02# => X"494e4700",
		16#4e03# => X"55736572",
		16#4e04# => X"5f54696d",
		16#4e05# => X"653a2025",
		16#4e06# => X"6c642c20",
		16#4e07# => X"54696d65",
		16#4e08# => X"2f52756e",
		16#4e09# => X"3a20256c",
		16#4e0a# => X"640a0000",
		16#4e0b# => X"4d696372",
		16#4e0c# => X"6f736563",
		16#4e0d# => X"6f6e6473",
		16#4e0e# => X"20666f72",
		16#4e0f# => X"206f6e65",
		16#4e10# => X"2072756e",
		16#4e11# => X"20746872",
		16#4e12# => X"6f756768",
		16#4e13# => X"20446872",
		16#4e14# => X"7973746f",
		16#4e15# => X"6e653a20",
		16#4e16# => X"256c640a",
		16#4e17# => X"00000000",
		16#4e18# => X"44687279",
		16#4e19# => X"73746f6e",
		16#4e1a# => X"65732070",
		16#4e1b# => X"65722053",
		16#4e1c# => X"65636f6e",
		16#4e1d# => X"643a2020",
		16#4e1e# => X"20202020",
		16#4e1f# => X"20202020",
		16#4e20# => X"20202020",
		16#4e21# => X"20202020",
		16#4e22# => X"20202020",
		16#4e23# => X"256c640a",
		16#4e24# => X"00000000",
		16#4e25# => X"44485259",
		16#4e26# => X"53544f4e",
		16#4e27# => X"45205052",
		16#4e28# => X"4f475241",
		16#4e29# => X"4d2c2031",
		16#4e2a# => X"27535420",
		16#4e2b# => X"53545249",
		16#4e2c# => X"4e470000",
		16#4e2d# => X"44485259",
		16#4e2e# => X"53544f4e",
		16#4e2f# => X"45205052",
		16#4e30# => X"4f475241",
		16#4e31# => X"4d2c2032",
		16#4e32# => X"274e4420",
		16#4e33# => X"53545249",
		16#4e34# => X"4e470000",
		16#4e35# => X"44485259",
		16#4e36# => X"53544f4e",
		16#4e37# => X"45205052",
		16#4e38# => X"4f475241",
		16#4e39# => X"4d2c2033",
		16#4e3a# => X"27524420",
		16#4e3b# => X"53545249",
		16#4e3c# => X"4e470000",
		16#4e3d# => X"494e4600",
		16#4e3e# => X"696e6600",
		16#4e3f# => X"4e414e00",
		16#4e40# => X"6e616e00",
		16#4e41# => X"30313233",
		16#4e42# => X"34353637",
		16#4e43# => X"38396162",
		16#4e44# => X"63646566",
		16#4e45# => X"00000000",
		16#4e46# => X"30313233",
		16#4e47# => X"34353637",
		16#4e48# => X"38394142",
		16#4e49# => X"43444546",
		16#4e4a# => X"00000000",
		16#4e4b# => X"30000000",
		16#4e4c# => X"204e614e",
		16#4e4d# => X"20000000",
		16#4e4e# => X"202d496e",
		16#4e4f# => X"66696e69",
		16#4e50# => X"74792000",
		16#4e51# => X"20496e66",
		16#4e52# => X"696e6974",
		16#4e53# => X"79200000",
		16#4e54# => X"4e614e00",
		16#4e55# => X"45256400",
		16#4e56# => X"43000000",
		16#4e57# => X"504f5349",
		16#4e58# => X"58000000",
		16#4e59# => X"2e000000",
		16#4e5a# => X"496d706c",
		16#4e5b# => X"656d656e",
		16#4e5c# => X"74206d61",
		16#4e5d# => X"696e2829",
		16#4e5e# => X"2c20666f",
		16#4e5f# => X"6f210000",
		16#4e60# => X"706e5f62",
		16#4e61# => X"6567696e",
		16#4e62# => X"5f706172",
		16#4e63# => X"616c6c65",
		16#4e64# => X"6c3a2045",
		16#4e65# => X"52524f52",
		16#4e66# => X"206e756d",
		16#4e67# => X"62657220",
		16#4e68# => X"6f662043",
		16#4e69# => X"6f505573",
		16#4e6a# => X"20656974",
		16#4e6b# => X"68657220",
		16#4e6c# => X"746f6f20",
		16#4e6d# => X"62696720",
		16#4e6e# => X"6f72206e",
		16#4e6f# => X"6f6e2070",
		16#4e70# => X"6c617573",
		16#4e71# => X"69626c65",
		16#4e72# => X"2076616c",
		16#4e73# => X"7565202d",
		16#4e74# => X"206e756d",
		16#4e75# => X"4350553a",
		16#4e76# => X"2025640d",
		16#4e77# => X"0a000000",
		16#4e78# => X"53746172",
		16#4e79# => X"74696e67",
		16#4e7a# => X"20436f50",
		16#4e7b# => X"55733a20",
		16#4e7c# => X"30782578",
		16#4e7d# => X"2c204a75",
		16#4e7e# => X"6d702061",
		16#4e7f# => X"64647265",
		16#4e80# => X"73733a20",
		16#4e81# => X"30782530",
		16#4e82# => X"38780d0a",
		16#4e83# => X"00000000",
		16#4e84# => X"706e5f62",
		16#4e85# => X"6567696e",
		16#4e86# => X"5f706172",
		16#4e87# => X"616c6c65",
		16#4e88# => X"6c3a2045",
		16#4e89# => X"52524f52",
		16#4e8a# => X"20636f75",
		16#4e8b# => X"6c64206e",
		16#4e8c# => X"6f742066",
		16#4e8d# => X"696e6420",
		16#4e8e# => X"656e6f75",
		16#4e8f# => X"67682043",
		16#4e90# => X"6f505573",
		16#4e91# => X"0d000000",
		16#4e92# => X"706e7468",
		16#4e93# => X"72656164",
		16#4e94# => X"5f637265",
		16#4e95# => X"6174653a",
		16#4e96# => X"20706e6d",
		16#4e97# => X"3263703a",
		16#4e98# => X"20307825",
		16#4e99# => X"782c2070",
		16#4e9a# => X"6e63656e",
		16#4e9b# => X"3a203078",
		16#4e9c# => X"25780d0a",
		16#4e9d# => X"00000000",
		16#4e9e# => X"706e7468",
		16#4e9f# => X"72656164",
		16#4ea0# => X"5f637265",
		16#4ea1# => X"6174653a",
		16#4ea2# => X"20537461",
		16#4ea3# => X"7274696e",
		16#4ea4# => X"67204350",
		16#4ea5# => X"5525642c",
		16#4ea6# => X"204a756d",
		16#4ea7# => X"70206164",
		16#4ea8# => X"64726573",
		16#4ea9# => X"73203078",
		16#4eaa# => X"25303878",
		16#4eab# => X"2c204172",
		16#4eac# => X"67206164",
		16#4ead# => X"64726573",
		16#4eae# => X"73203078",
		16#4eaf# => X"25303878",
		16#4eb0# => X"0d0a0000",
		16#4eb1# => X"706e7468",
		16#4eb2# => X"72656164",
		16#4eb3# => X"5f637265",
		16#4eb4# => X"6174653a",
		16#4eb5# => X"20746872",
		16#4eb6# => X"6561645f",
		16#4eb7# => X"726f7574",
		16#4eb8# => X"696e6520",
		16#4eb9# => X"30782530",
		16#4eba# => X"38782c20",
		16#4ebb# => X"74687265",
		16#4ebc# => X"61645f61",
		16#4ebd# => X"72672030",
		16#4ebe# => X"78253038",
		16#4ebf# => X"780d0a00",
		16#4ec0# => X"706e7468",
		16#4ec1# => X"72656164",
		16#4ec2# => X"5f637265",
		16#4ec3# => X"6174653a",
		16#4ec4# => X"20537461",
		16#4ec5# => X"7274696e",
		16#4ec6# => X"67204365",
		16#4ec7# => X"50553a20",
		16#4ec8# => X"4a756d70",
		16#4ec9# => X"20616464",
		16#4eca# => X"72657373",
		16#4ecb# => X"20307825",
		16#4ecc# => X"3038780d",
		16#4ecd# => X"0a000000",
		16#4ece# => X"48656170",
		16#4ecf# => X"20616e64",
		16#4ed0# => X"20737461",
		16#4ed1# => X"636b2063",
		16#4ed2# => X"6f6c6c69",
		16#4ed3# => X"73696f6e",
		16#4ed4# => X"00000000",
		16#4ed5# => X"00000000",
		16#4ed6# => X"641b0010",
		16#4ed7# => X"e42c0010",
		16#4ed8# => X"e42c0010",
		16#4ed9# => X"781b0010",
		16#4eda# => X"e42c0010",
		16#4edb# => X"e42c0010",
		16#4edc# => X"e42c0010",
		16#4edd# => X"181b0010",
		16#4ede# => X"e42c0010",
		16#4edf# => X"e42c0010",
		16#4ee0# => X"801b0010",
		16#4ee1# => X"a01b0010",
		16#4ee2# => X"e42c0010",
		16#4ee3# => X"981b0010",
		16#4ee4# => X"a81b0010",
		16#4ee5# => X"e42c0010",
		16#4ee6# => X"141c0010",
		16#4ee7# => X"1c1c0010",
		16#4ee8# => X"1c1c0010",
		16#4ee9# => X"1c1c0010",
		16#4eea# => X"1c1c0010",
		16#4eeb# => X"1c1c0010",
		16#4eec# => X"1c1c0010",
		16#4eed# => X"1c1c0010",
		16#4eee# => X"1c1c0010",
		16#4eef# => X"1c1c0010",
		16#4ef0# => X"e42c0010",
		16#4ef1# => X"e42c0010",
		16#4ef2# => X"e42c0010",
		16#4ef3# => X"e42c0010",
		16#4ef4# => X"e42c0010",
		16#4ef5# => X"e42c0010",
		16#4ef6# => X"e42c0010",
		16#4ef7# => X"28200010",
		16#4ef8# => X"e42c0010",
		16#4ef9# => X"b81c0010",
		16#4efa# => X"7c1f0010",
		16#4efb# => X"28200010",
		16#4efc# => X"28200010",
		16#4efd# => X"28200010",
		16#4efe# => X"e42c0010",
		16#4eff# => X"e42c0010",
		16#4f00# => X"e42c0010",
		16#4f01# => X"e42c0010",
		16#4f02# => X"581c0010",
		16#4f03# => X"e42c0010",
		16#4f04# => X"e42c0010",
		16#4f05# => X"88290010",
		16#4f06# => X"e42c0010",
		16#4f07# => X"e42c0010",
		16#4f08# => X"e42c0010",
		16#4f09# => X"582a0010",
		16#4f0a# => X"e42c0010",
		16#4f0b# => X"a42a0010",
		16#4f0c# => X"e42c0010",
		16#4f0d# => X"e42c0010",
		16#4f0e# => X"b81a0010",
		16#4f0f# => X"e42c0010",
		16#4f10# => X"e42c0010",
		16#4f11# => X"e42c0010",
		16#4f12# => X"e42c0010",
		16#4f13# => X"e42c0010",
		16#4f14# => X"e42c0010",
		16#4f15# => X"e42c0010",
		16#4f16# => X"e42c0010",
		16#4f17# => X"28200010",
		16#4f18# => X"e42c0010",
		16#4f19# => X"b81c0010",
		16#4f1a# => X"801f0010",
		16#4f1b# => X"28200010",
		16#4f1c# => X"28200010",
		16#4f1d# => X"28200010",
		16#4f1e# => X"601c0010",
		16#4f1f# => X"801f0010",
		16#4f20# => X"a81c0010",
		16#4f21# => X"e42c0010",
		16#4f22# => X"8c1c0010",
		16#4f23# => X"e42c0010",
		16#4f24# => X"1c290010",
		16#4f25# => X"8c290010",
		16#4f26# => X"1c2a0010",
		16#4f27# => X"a81c0010",
		16#4f28# => X"e42c0010",
		16#4f29# => X"582a0010",
		16#4f2a# => X"741a0010",
		16#4f2b# => X"a82a0010",
		16#4f2c# => X"e42c0010",
		16#4f2d# => X"e42c0010",
		16#4f2e# => X"0c2b0010",
		16#4f2f# => X"e42c0010",
		16#4f30# => X"741a0010",
		16#4f31# => X"20202020",
		16#4f32# => X"20202020",
		16#4f33# => X"20202020",
		16#4f34# => X"20202020",
		16#4f35# => X"30303030",
		16#4f36# => X"30303030",
		16#4f37# => X"30303030",
		16#4f38# => X"30303030",
		16#4f39# => X"00000000",
		16#4f3a# => X"00000000",
		16#4f3b# => X"00000000",
		16#4f3c# => X"00000000",
		16#4f3d# => X"00000000",
		16#4f3e# => X"00000000",
		16#4f3f# => X"00000000",
		16#4f40# => X"00000000",
		16#4f41# => X"00000000",
		16#4f42# => X"0080ff3f",
		16#4f43# => X"7665924a",
		16#4f44# => X"4a803f15",
		16#4f45# => X"4cc99a97",
		16#4f46# => X"208a0252",
		16#4f47# => X"60c42575",
		16#4f48# => X"326a52ce",
		16#4f49# => X"9a32ce28",
		16#4f4a# => X"4da7e45d",
		16#4f4b# => X"3dc55d3b",
		16#4f4c# => X"8b9e925a",
		16#4f4d# => X"6c52ce50",
		16#4f4e# => X"8bf1283d",
		16#4f4f# => X"0d65170c",
		16#4f50# => X"75818675",
		16#4f51# => X"76c9484d",
		16#4f52# => X"669cf858",
		16#4f53# => X"50bc545c",
		16#4f54# => X"65ccc691",
		16#4f55# => X"0ea6aea0",
		16#4f56# => X"19e3a346",
		16#4f57# => X"1e85b7ea",
		16#4f58# => X"fe981b90",
		16#4f59# => X"bbdd8dde",
		16#4f5a# => X"f99dfbeb",
		16#4f5b# => X"7eaa5143",
		16#4f5c# => X"35023701",
		16#4f5d# => X"b1366c33",
		16#4f5e# => X"6fc6df8c",
		16#4f5f# => X"e980c947",
		16#4f60# => X"ba93a841",
		16#4f61# => X"f850fb25",
		16#4f62# => X"6bc7716b",
		16#4f63# => X"bf3cd5a6",
		16#4f64# => X"cfff491f",
		16#4f65# => X"78c2d340",
		16#4f66# => X"00000000",
		16#4f67# => X"00000000",
		16#4f68# => X"20f09db5",
		16#4f69# => X"702ba8ad",
		16#4f6a# => X"c59d6940",
		16#4f6b# => X"00000000",
		16#4f6c# => X"00000000",
		16#4f6d# => X"00000000",
		16#4f6e# => X"0004bfc9",
		16#4f6f# => X"1b8e3440",
		16#4f70# => X"00000000",
		16#4f71# => X"00000000",
		16#4f72# => X"00000000",
		16#4f73# => X"00000020",
		16#4f74# => X"bcbe1940",
		16#4f75# => X"00000000",
		16#4f76# => X"00000000",
		16#4f77# => X"00000000",
		16#4f78# => X"00000000",
		16#4f79# => X"409c0c40",
		16#4f7a# => X"00000000",
		16#4f7b# => X"00000000",
		16#4f7c# => X"00000000",
		16#4f7d# => X"00000000",
		16#4f7e# => X"00c80540",
		16#4f7f# => X"00000000",
		16#4f80# => X"00000000",
		16#4f81# => X"00000000",
		16#4f82# => X"00000000",
		16#4f83# => X"00a00240",
		16#4f84# => X"fffffeff",
		16#4f85# => X"fcfff8ff",
		16#4f86# => X"f0ffe0ff",
		16#4f87# => X"c0ff80ff",
		16#4f88# => X"00ff00fe",
		16#4f89# => X"00fc00f8",
		16#4f8a# => X"00f000e0",
		16#4f8b# => X"00c00080",
		16#4f8c# => X"00000000",
		16#4f8d# => X"3020fccf",
		16#4f8e# => X"c3a12381",
		16#4f8f# => X"e32dde9f",
		16#4f90# => X"ced2c804",
		16#4f91# => X"dda6d80a",
		16#4f92# => X"6482cbd2",
		16#4f93# => X"eaf2d412",
		16#4f94# => X"2549e42d",
		16#4f95# => X"36344f53",
		16#4f96# => X"aece6b25",
		16#4f97# => X"3ff598f6",
		16#4f98# => X"d36b5801",
		16#4f99# => X"a687bdc0",
		16#4f9a# => X"57daa582",
		16#4f9b# => X"a6a2b532",
		16#4f9c# => X"31e7d404",
		16#4f9d# => X"f2e332d3",
		16#4f9e# => X"32711cd2",
		16#4f9f# => X"23db32ee",
		16#4fa0# => X"49905a39",
		16#4fa1# => X"3ea20853",
		16#4fa2# => X"fbfe5511",
		16#4fa3# => X"91fa3919",
		16#4fa4# => X"7a632543",
		16#4fa5# => X"31c0ac3c",
		16#4fa6# => X"6de2dedb",
		16#4fa7# => X"5dd0f6b3",
		16#4fa8# => X"7caca0e4",
		16#4fa9# => X"bc647c46",
		16#4faa# => X"d0dd553e",
		16#4fab# => X"202a2462",
		16#4fac# => X"b347d798",
		16#4fad# => X"233fa5e9",
		16#4fae# => X"39a527ea",
		16#4faf# => X"7fa82a3f",
		16#4fb0# => X"5b0bf24a",
		16#4fb1# => X"81a5ed18",
		16#4fb2# => X"de67ba94",
		16#4fb3# => X"3945ad1e",
		16#4fb4# => X"b1cf943f",
		16#4fb5# => X"71bfb3a9",
		16#4fb6# => X"897968be",
		16#4fb7# => X"2e4c5be1",
		16#4fb8# => X"4dc4be94",
		16#4fb9# => X"95e6c93f",
		16#4fba# => X"4d3d3d7c",
		16#4fbb# => X"ba362b0d",
		16#4fbc# => X"c2fdfcce",
		16#4fbd# => X"61841177",
		16#4fbe# => X"ccabe43f",
		16#4fbf# => X"55c1a8a4",
		16#4fc0# => X"4e401361",
		16#4fc1# => X"c3d32b65",
		16#4fc2# => X"19e25817",
		16#4fc3# => X"b7d1f13f",
		16#4fc4# => X"0ad7a370",
		16#4fc5# => X"3d0ad7a3",
		16#4fc6# => X"703d0ad7",
		16#4fc7# => X"a3703d0a",
		16#4fc8# => X"d7a3f83f",
		16#4fc9# => X"cdcccccc",
		16#4fca# => X"cccccccc",
		16#4fcb# => X"cccccccc",
		16#4fcc# => X"cccccccc",
		16#4fcd# => X"ccccfb3f",
		16#4fce# => X"05000000",
		16#4fcf# => X"19000000",
		16#4fd0# => X"7d000000",
		16#4fd1# => X"00000000",
		16#4fd2# => X"00000000",
		16#4fd3# => X"0000f03f",
		16#4fd4# => X"00000000",
		16#4fd5# => X"00002440",
		16#4fd6# => X"00000000",
		16#4fd7# => X"00005940",
		16#4fd8# => X"00000000",
		16#4fd9# => X"00408f40",
		16#4fda# => X"00000000",
		16#4fdb# => X"0088c340",
		16#4fdc# => X"00000000",
		16#4fdd# => X"006af840",
		16#4fde# => X"00000000",
		16#4fdf# => X"80842e41",
		16#4fe0# => X"00000000",
		16#4fe1# => X"d0126341",
		16#4fe2# => X"00000000",
		16#4fe3# => X"84d79741",
		16#4fe4# => X"00000000",
		16#4fe5# => X"65cdcd41",
		16#4fe6# => X"00000020",
		16#4fe7# => X"5fa00242",
		16#4fe8# => X"000000e8",
		16#4fe9# => X"76483742",
		16#4fea# => X"000000a2",
		16#4feb# => X"941a6d42",
		16#4fec# => X"000040e5",
		16#4fed# => X"9c30a242",
		16#4fee# => X"0000901e",
		16#4fef# => X"c4bcd642",
		16#4ff0# => X"00003426",
		16#4ff1# => X"f56b0c43",
		16#4ff2# => X"0080e037",
		16#4ff3# => X"79c34143",
		16#4ff4# => X"00a0d885",
		16#4ff5# => X"57347643",
		16#4ff6# => X"00c84e67",
		16#4ff7# => X"6dc1ab43",
		16#4ff8# => X"003d9160",
		16#4ff9# => X"e458e143",
		16#4ffa# => X"408cb578",
		16#4ffb# => X"1daf1544",
		16#4ffc# => X"50efe2d6",
		16#4ffd# => X"e41a4b44",
		16#4ffe# => X"92d54d06",
		16#4fff# => X"cff08044",
		16#5000# => X"f64ae1c7",
		16#5001# => X"022db544",
		16#5002# => X"b49dd979",
		16#5003# => X"4378ea44",
		16#5004# => X"bc89d897",
		16#5005# => X"b2d29c3c",
		16#5006# => X"33a7a8d5",
		16#5007# => X"23f64939",
		16#5008# => X"3da7f444",
		16#5009# => X"fd0fa532",
		16#500a# => X"9d978ccf",
		16#500b# => X"08ba5b25",
		16#500c# => X"436fac64",
		16#500d# => X"2806c80a",
		16#500e# => X"0080e037",
		16#500f# => X"79c34143",
		16#5010# => X"176e05b5",
		16#5011# => X"b5b89346",
		16#5012# => X"f5f93fe9",
		16#5013# => X"034f384d",
		16#5014# => X"321d30f9",
		16#5015# => X"4877825a",
		16#5016# => X"3cbf737f",
		16#5017# => X"dd4f1575",
		16#5018# => X"80900010",
		16#5019# => X"3ca20010",
		16#501a# => X"3ca20010",
		16#501b# => X"94900010",
		16#501c# => X"3ca20010",
		16#501d# => X"3ca20010",
		16#501e# => X"3ca20010",
		16#501f# => X"34900010",
		16#5020# => X"3ca20010",
		16#5021# => X"3ca20010",
		16#5022# => X"9c900010",
		16#5023# => X"bc900010",
		16#5024# => X"3ca20010",
		16#5025# => X"b4900010",
		16#5026# => X"c4900010",
		16#5027# => X"3ca20010",
		16#5028# => X"30910010",
		16#5029# => X"38910010",
		16#502a# => X"38910010",
		16#502b# => X"38910010",
		16#502c# => X"38910010",
		16#502d# => X"38910010",
		16#502e# => X"38910010",
		16#502f# => X"38910010",
		16#5030# => X"38910010",
		16#5031# => X"38910010",
		16#5032# => X"3ca20010",
		16#5033# => X"3ca20010",
		16#5034# => X"3ca20010",
		16#5035# => X"3ca20010",
		16#5036# => X"3ca20010",
		16#5037# => X"3ca20010",
		16#5038# => X"3ca20010",
		16#5039# => X"44950010",
		16#503a# => X"3ca20010",
		16#503b# => X"d4910010",
		16#503c# => X"98940010",
		16#503d# => X"44950010",
		16#503e# => X"44950010",
		16#503f# => X"44950010",
		16#5040# => X"3ca20010",
		16#5041# => X"3ca20010",
		16#5042# => X"3ca20010",
		16#5043# => X"3ca20010",
		16#5044# => X"74910010",
		16#5045# => X"3ca20010",
		16#5046# => X"3ca20010",
		16#5047# => X"e09e0010",
		16#5048# => X"3ca20010",
		16#5049# => X"3ca20010",
		16#504a# => X"3ca20010",
		16#504b# => X"b09f0010",
		16#504c# => X"3ca20010",
		16#504d# => X"fc9f0010",
		16#504e# => X"3ca20010",
		16#504f# => X"3ca20010",
		16#5050# => X"d48f0010",
		16#5051# => X"3ca20010",
		16#5052# => X"3ca20010",
		16#5053# => X"3ca20010",
		16#5054# => X"3ca20010",
		16#5055# => X"3ca20010",
		16#5056# => X"3ca20010",
		16#5057# => X"3ca20010",
		16#5058# => X"3ca20010",
		16#5059# => X"44950010",
		16#505a# => X"3ca20010",
		16#505b# => X"d4910010",
		16#505c# => X"9c940010",
		16#505d# => X"44950010",
		16#505e# => X"44950010",
		16#505f# => X"44950010",
		16#5060# => X"7c910010",
		16#5061# => X"9c940010",
		16#5062# => X"c4910010",
		16#5063# => X"3ca20010",
		16#5064# => X"a8910010",
		16#5065# => X"3ca20010",
		16#5066# => X"749e0010",
		16#5067# => X"e49e0010",
		16#5068# => X"749f0010",
		16#5069# => X"c4910010",
		16#506a# => X"3ca20010",
		16#506b# => X"b09f0010",
		16#506c# => X"908f0010",
		16#506d# => X"00a00010",
		16#506e# => X"3ca20010",
		16#506f# => X"3ca20010",
		16#5070# => X"64a00010",
		16#5071# => X"3ca20010",
		16#5072# => X"908f0010",
		16#5073# => X"20202020",
		16#5074# => X"20202020",
		16#5075# => X"20202020",
		16#5076# => X"20202020",
		16#5077# => X"30303030",
		16#5078# => X"30303030",
		16#5079# => X"30303030",
		16#507a# => X"30303030",
		16#507b# => X"14b10010",
		16#507c# => X"18b90010",
		16#507d# => X"18b90010",
		16#507e# => X"28b10010",
		16#507f# => X"18b90010",
		16#5080# => X"18b90010",
		16#5081# => X"18b90010",
		16#5082# => X"c8b00010",
		16#5083# => X"18b90010",
		16#5084# => X"18b90010",
		16#5085# => X"30b10010",
		16#5086# => X"48b10010",
		16#5087# => X"18b90010",
		16#5088# => X"40b10010",
		16#5089# => X"50b10010",
		16#508a# => X"18b90010",
		16#508b# => X"acb10010",
		16#508c# => X"b4b10010",
		16#508d# => X"b4b10010",
		16#508e# => X"b4b10010",
		16#508f# => X"b4b10010",
		16#5090# => X"b4b10010",
		16#5091# => X"b4b10010",
		16#5092# => X"b4b10010",
		16#5093# => X"b4b10010",
		16#5094# => X"b4b10010",
		16#5095# => X"18b90010",
		16#5096# => X"18b90010",
		16#5097# => X"18b90010",
		16#5098# => X"18b90010",
		16#5099# => X"18b90010",
		16#509a# => X"18b90010",
		16#509b# => X"18b90010",
		16#509c# => X"18b90010",
		16#509d# => X"18b90010",
		16#509e# => X"24b20010",
		16#509f# => X"44b20010",
		16#50a0# => X"18b90010",
		16#50a1# => X"18b90010",
		16#50a2# => X"18b90010",
		16#50a3# => X"18b90010",
		16#50a4# => X"18b90010",
		16#50a5# => X"18b90010",
		16#50a6# => X"18b90010",
		16#50a7# => X"18b90010",
		16#50a8# => X"18b90010",
		16#50a9# => X"18b90010",
		16#50aa# => X"48b30010",
		16#50ab# => X"18b90010",
		16#50ac# => X"18b90010",
		16#50ad# => X"18b90010",
		16#50ae# => X"04b40010",
		16#50af# => X"18b90010",
		16#50b0# => X"d8b60010",
		16#50b1# => X"18b90010",
		16#50b2# => X"18b90010",
		16#50b3# => X"78b00010",
		16#50b4# => X"18b90010",
		16#50b5# => X"18b90010",
		16#50b6# => X"18b90010",
		16#50b7# => X"18b90010",
		16#50b8# => X"18b90010",
		16#50b9# => X"18b90010",
		16#50ba# => X"18b90010",
		16#50bb# => X"18b90010",
		16#50bc# => X"18b90010",
		16#50bd# => X"18b90010",
		16#50be# => X"24b20010",
		16#50bf# => X"48b20010",
		16#50c0# => X"18b90010",
		16#50c1# => X"18b90010",
		16#50c2# => X"18b90010",
		16#50c3# => X"e4b10010",
		16#50c4# => X"48b20010",
		16#50c5# => X"14b20010",
		16#50c6# => X"18b90010",
		16#50c7# => X"04b20010",
		16#50c8# => X"18b90010",
		16#50c9# => X"e8b20010",
		16#50ca# => X"4cb30010",
		16#50cb# => X"d4b30010",
		16#50cc# => X"14b20010",
		16#50cd# => X"18b90010",
		16#50ce# => X"04b40010",
		16#50cf# => X"4cb00010",
		16#50d0# => X"dcb60010",
		16#50d1# => X"18b90010",
		16#50d2# => X"18b90010",
		16#50d3# => X"38b70010",
		16#50d4# => X"18b90010",
		16#50d5# => X"4cb00010",
		16#50d6# => X"20202020",
		16#50d7# => X"20202020",
		16#50d8# => X"20202020",
		16#50d9# => X"20202020",
		16#50da# => X"30303030",
		16#50db# => X"30303030",
		16#50dc# => X"30303030",
		16#50dd# => X"30303030",
		16#50de# => X"00202020",
		16#50df# => X"20202020",
		16#50e0# => X"20202828",
		16#50e1# => X"28282820",
		16#50e2# => X"20202020",
		16#50e3# => X"20202020",
		16#50e4# => X"20202020",
		16#50e5# => X"20202020",
		16#50e6# => X"20881010",
		16#50e7# => X"10101010",
		16#50e8# => X"10101010",
		16#50e9# => X"10101010",
		16#50ea# => X"10040404",
		16#50eb# => X"04040404",
		16#50ec# => X"04040410",
		16#50ed# => X"10101010",
		16#50ee# => X"10104141",
		16#50ef# => X"41414141",
		16#50f0# => X"01010101",
		16#50f1# => X"01010101",
		16#50f2# => X"01010101",
		16#50f3# => X"01010101",
		16#50f4# => X"01010101",
		16#50f5# => X"10101010",
		16#50f6# => X"10104242",
		16#50f7# => X"42424242",
		16#50f8# => X"02020202",
		16#50f9# => X"02020202",
		16#50fa# => X"02020202",
		16#50fb# => X"02020202",
		16#50fc# => X"02020202",
		16#50fd# => X"10101010",
		16#50fe# => X"20000000",
		16#50ff# => X"00000000",
		16#5100# => X"00000000",
		16#5101# => X"00000000",
		16#5102# => X"00000000",
		16#5103# => X"00000000",
		16#5104# => X"00000000",
		16#5105# => X"00000000",
		16#5106# => X"00000000",
		16#5107# => X"00000000",
		16#5108# => X"00000000",
		16#5109# => X"00000000",
		16#510a# => X"00000000",
		16#510b# => X"00000000",
		16#510c# => X"00000000",
		16#510d# => X"00000000",
		16#510e# => X"00000000",
		16#510f# => X"00000000",
		16#5110# => X"00000000",
		16#5111# => X"00000000",
		16#5112# => X"00000000",
		16#5113# => X"00000000",
		16#5114# => X"00000000",
		16#5115# => X"00000000",
		16#5116# => X"00000000",
		16#5117# => X"00000000",
		16#5118# => X"00000000",
		16#5119# => X"00000000",
		16#511a# => X"00000000",
		16#511b# => X"00000000",
		16#511c# => X"00000000",
		16#511d# => X"00000000",
		16#511e# => X"00000000",
		16#511f# => X"2cc60010",
		16#5120# => X"30ce0010",
		16#5121# => X"30ce0010",
		16#5122# => X"40c60010",
		16#5123# => X"30ce0010",
		16#5124# => X"30ce0010",
		16#5125# => X"30ce0010",
		16#5126# => X"e0c50010",
		16#5127# => X"30ce0010",
		16#5128# => X"30ce0010",
		16#5129# => X"48c60010",
		16#512a# => X"60c60010",
		16#512b# => X"30ce0010",
		16#512c# => X"58c60010",
		16#512d# => X"68c60010",
		16#512e# => X"30ce0010",
		16#512f# => X"c4c60010",
		16#5130# => X"ccc60010",
		16#5131# => X"ccc60010",
		16#5132# => X"ccc60010",
		16#5133# => X"ccc60010",
		16#5134# => X"ccc60010",
		16#5135# => X"ccc60010",
		16#5136# => X"ccc60010",
		16#5137# => X"ccc60010",
		16#5138# => X"ccc60010",
		16#5139# => X"30ce0010",
		16#513a# => X"30ce0010",
		16#513b# => X"30ce0010",
		16#513c# => X"30ce0010",
		16#513d# => X"30ce0010",
		16#513e# => X"30ce0010",
		16#513f# => X"30ce0010",
		16#5140# => X"30ce0010",
		16#5141# => X"30ce0010",
		16#5142# => X"3cc70010",
		16#5143# => X"5cc70010",
		16#5144# => X"30ce0010",
		16#5145# => X"30ce0010",
		16#5146# => X"30ce0010",
		16#5147# => X"30ce0010",
		16#5148# => X"30ce0010",
		16#5149# => X"30ce0010",
		16#514a# => X"30ce0010",
		16#514b# => X"30ce0010",
		16#514c# => X"30ce0010",
		16#514d# => X"30ce0010",
		16#514e# => X"60c80010",
		16#514f# => X"30ce0010",
		16#5150# => X"30ce0010",
		16#5151# => X"30ce0010",
		16#5152# => X"1cc90010",
		16#5153# => X"30ce0010",
		16#5154# => X"f0cb0010",
		16#5155# => X"30ce0010",
		16#5156# => X"30ce0010",
		16#5157# => X"90c50010",
		16#5158# => X"30ce0010",
		16#5159# => X"30ce0010",
		16#515a# => X"30ce0010",
		16#515b# => X"30ce0010",
		16#515c# => X"30ce0010",
		16#515d# => X"30ce0010",
		16#515e# => X"30ce0010",
		16#515f# => X"30ce0010",
		16#5160# => X"30ce0010",
		16#5161# => X"30ce0010",
		16#5162# => X"3cc70010",
		16#5163# => X"60c70010",
		16#5164# => X"30ce0010",
		16#5165# => X"30ce0010",
		16#5166# => X"30ce0010",
		16#5167# => X"fcc60010",
		16#5168# => X"60c70010",
		16#5169# => X"2cc70010",
		16#516a# => X"30ce0010",
		16#516b# => X"1cc70010",
		16#516c# => X"30ce0010",
		16#516d# => X"00c80010",
		16#516e# => X"64c80010",
		16#516f# => X"ecc80010",
		16#5170# => X"2cc70010",
		16#5171# => X"30ce0010",
		16#5172# => X"1cc90010",
		16#5173# => X"64c50010",
		16#5174# => X"f4cb0010",
		16#5175# => X"30ce0010",
		16#5176# => X"30ce0010",
		16#5177# => X"50cc0010",
		16#5178# => X"30ce0010",
		16#5179# => X"64c50010",
		16#517a# => X"20202020",
		16#517b# => X"20202020",
		16#517c# => X"20202020",
		16#517d# => X"20202020",
		16#517e# => X"30303030",
		16#517f# => X"30303030",
		16#5180# => X"30303030",
		16#5181# => X"30303030",
		16#5182# => X"ace90010",
		16#5183# => X"c0e80010",
		16#5184# => X"cce80010",
		16#5185# => X"c0e80010",
		16#5186# => X"98e90010",
		16#5187# => X"c0e80010",
		16#5188# => X"cce80010",
		16#5189# => X"ace90010",
		16#518a# => X"ace90010",
		16#518b# => X"98e90010",
		16#518c# => X"cce80010",
		16#518d# => X"98e80010",
		16#518e# => X"98e80010",
		16#518f# => X"98e80010",
		16#5190# => X"d4e80010",
		16#5191# => X"a0ef0010",
		16#5192# => X"a0ef0010",
		16#5193# => X"c4ef0010",
		16#5194# => X"94ef0010",
		16#5195# => X"94ef0010",
		16#5196# => X"84f00010",
		16#5197# => X"c4ef0010",
		16#5198# => X"94ef0010",
		16#5199# => X"84f00010",
		16#519a# => X"94ef0010",
		16#519b# => X"c4ef0010",
		16#519c# => X"90ef0010",
		16#519d# => X"90ef0010",
		16#519e# => X"90ef0010",
		16#519f# => X"84f00010",
		16#51a0# => X"10060110",
		16#51a1# => X"10060110",
		16#51a2# => X"0c060110",
		16#51a3# => X"c0050110",
		16#51a4# => X"c0050110",
		16#51a5# => X"80080110",
		16#51a6# => X"0c060110",
		16#51a7# => X"c0050110",
		16#51a8# => X"80080110",
		16#51a9# => X"c0050110",
		16#51aa# => X"0c060110",
		16#51ab# => X"bc050110",
		16#51ac# => X"bc050110",
		16#51ad# => X"bc050110",
		16#51ae# => X"80080110",
		16#51af# => X"00010202",
		16#51b0# => X"03030303",
		16#51b1# => X"04040404",
		16#51b2# => X"04040404",
		16#51b3# => X"05050505",
		16#51b4# => X"05050505",
		16#51b5# => X"05050505",
		16#51b6# => X"05050505",
		16#51b7# => X"06060606",
		16#51b8# => X"06060606",
		16#51b9# => X"06060606",
		16#51ba# => X"06060606",
		16#51bb# => X"06060606",
		16#51bc# => X"06060606",
		16#51bd# => X"06060606",
		16#51be# => X"06060606",
		16#51bf# => X"07070707",
		16#51c0# => X"07070707",
		16#51c1# => X"07070707",
		16#51c2# => X"07070707",
		16#51c3# => X"07070707",
		16#51c4# => X"07070707",
		16#51c5# => X"07070707",
		16#51c6# => X"07070707",
		16#51c7# => X"07070707",
		16#51c8# => X"07070707",
		16#51c9# => X"07070707",
		16#51ca# => X"07070707",
		16#51cb# => X"07070707",
		16#51cc# => X"07070707",
		16#51cd# => X"07070707",
		16#51ce# => X"07070707",
		16#51cf# => X"08080808",
		16#51d0# => X"08080808",
		16#51d1# => X"08080808",
		16#51d2# => X"08080808",
		16#51d3# => X"08080808",
		16#51d4# => X"08080808",
		16#51d5# => X"08080808",
		16#51d6# => X"08080808",
		16#51d7# => X"08080808",
		16#51d8# => X"08080808",
		16#51d9# => X"08080808",
		16#51da# => X"08080808",
		16#51db# => X"08080808",
		16#51dc# => X"08080808",
		16#51dd# => X"08080808",
		16#51de# => X"08080808",
		16#51df# => X"08080808",
		16#51e0# => X"08080808",
		16#51e1# => X"08080808",
		16#51e2# => X"08080808",
		16#51e3# => X"08080808",
		16#51e4# => X"08080808",
		16#51e5# => X"08080808",
		16#51e6# => X"08080808",
		16#51e7# => X"08080808",
		16#51e8# => X"08080808",
		16#51e9# => X"08080808",
		16#51ea# => X"08080808",
		16#51eb# => X"08080808",
		16#51ec# => X"08080808",
		16#51ed# => X"08080808",
		16#51ee# => X"08080808",
		16#51ef# => X"10000000",
		16#51f0# => X"00000000",
		16#51f1# => X"017a5200",
		16#51f2# => X"017c0101",
		16#51f3# => X"1b0d0200",
		16#51f4# => X"4c000000",
		16#51f5# => X"18000000",
		16#51f6# => X"0c8fffff",
		16#51f7# => X"dc050000",
		16#51f8# => X"00440e30",
		16#51f9# => X"70960897",
		16#51fa# => X"09810188",
		16#51fb# => X"02890392",
		16#51fc# => X"04930594",
		16#51fd# => X"06950798",
		16#51fe# => X"0a990b9a",
		16#51ff# => X"0c037002",
		16#5200# => X"0ac144c8",
		16#5201# => X"44c944d2",
		16#5202# => X"44d344d4",
		16#5203# => X"44d544d6",
		16#5204# => X"44d744d8",
		16#5205# => X"44d944da",
		16#5206# => X"440e0044",
		16#5207# => X"0b000000",
		16#5208# => X"50000000",
		16#5209# => X"68000000",
		16#520a# => X"9894ffff",
		16#520b# => X"00050000",
		16#520c# => X"00440e50",
		16#520d# => X"74880289",
		16#520e# => X"03930599",
		16#520f# => X"0b810192",
		16#5210# => X"04940695",
		16#5211# => X"07960897",
		16#5212# => X"09980a9a",
		16#5213# => X"0c9b0d03",
		16#5214# => X"20010ac1",
		16#5215# => X"44c844c9",
		16#5216# => X"44d244d3",
		16#5217# => X"44d444d5",
		16#5218# => X"44d644d7",
		16#5219# => X"44d844d9",
		16#521a# => X"44da44db",
		16#521b# => X"440e0044",
		16#521c# => X"0b000000",
		16#521d# => X"00000000",
		16#521e# => X"00000000",
		16#521f# => X"644b0110",
		16#5220# => X"cc4b0110",
		16#5221# => X"344c0110",
		16#5222# => X"00000000",
		16#5223# => X"00000000",
		16#5224# => X"00000000",
		16#5225# => X"00000000",
		16#5226# => X"00000000",
		16#5227# => X"00000000",
		16#5228# => X"00000000",
		16#5229# => X"00000000",
		16#522a# => X"00000000",
		16#522b# => X"00000000",
		16#522c# => X"00000000",
		16#522d# => X"00000000",
		16#522e# => X"00000000",
		16#522f# => X"00000000",
		16#5230# => X"00000000",
		16#5231# => X"00000000",
		16#5232# => X"00000000",
		16#5233# => X"00000000",
		16#5234# => X"00000000",
		16#5235# => X"00000000",
		16#5236# => X"00000000",
		16#5237# => X"00000000",
		16#5238# => X"00000000",
		16#5239# => X"00000000",
		16#523a# => X"00000000",
		16#523b# => X"00000000",
		16#523c# => X"00000000",
		16#523d# => X"00000000",
		16#523e# => X"00000000",
		16#523f# => X"00000000",
		16#5240# => X"00000000",
		16#5241# => X"00000000",
		16#5242# => X"00000000",
		16#5243# => X"00000000",
		16#5244# => X"00000000",
		16#5245# => X"00000000",
		16#5246# => X"00000000",
		16#5247# => X"00000000",
		16#5248# => X"01000000",
		16#5249# => X"00000000",
		16#524a# => X"0e33cdab",
		16#524b# => X"34126de6",
		16#524c# => X"ecde0500",
		16#524d# => X"0b000000",
		16#524e# => X"00000000",
		16#524f# => X"00000000",
		16#5250# => X"00000000",
		16#5251# => X"00000000",
		16#5252# => X"00000000",
		16#5253# => X"00000000",
		16#5254# => X"00000000",
		16#5255# => X"00000000",
		16#5256# => X"00000000",
		16#5257# => X"00000000",
		16#5258# => X"00000000",
		16#5259# => X"00000000",
		16#525a# => X"00000000",
		16#525b# => X"00000000",
		16#525c# => X"00000000",
		16#525d# => X"00000000",
		16#525e# => X"00000000",
		16#525f# => X"00000000",
		16#5260# => X"00000000",
		16#5261# => X"00000000",
		16#5262# => X"00000000",
		16#5263# => X"00000000",
		16#5264# => X"00000000",
		16#5265# => X"00000000",
		16#5266# => X"00000000",
		16#5267# => X"00000000",
		16#5268# => X"00000000",
		16#5269# => X"00000000",
		16#526a# => X"00000000",
		16#526b# => X"00000000",
		16#526c# => X"00000000",
		16#526d# => X"00000000",
		16#526e# => X"00000000",
		16#526f# => X"00000000",
		16#5270# => X"00000000",
		16#5271# => X"00000000",
		16#5272# => X"00000000",
		16#5273# => X"00000000",
		16#5274# => X"00000000",
		16#5275# => X"00000000",
		16#5276# => X"00000000",
		16#5277# => X"00000000",
		16#5278# => X"00000000",
		16#5279# => X"00000000",
		16#527a# => X"00000000",
		16#527b# => X"00000000",
		16#527c# => X"00000000",
		16#527d# => X"00000000",
		16#527e# => X"00000000",
		16#527f# => X"00000000",
		16#5280# => X"00000000",
		16#5281# => X"00000000",
		16#5282# => X"00000000",
		16#5283# => X"00000000",
		16#5284# => X"00000000",
		16#5285# => X"00000000",
		16#5286# => X"00000000",
		16#5287# => X"00000000",
		16#5288# => X"00000000",
		16#5289# => X"00000000",
		16#528a# => X"00000000",
		16#528b# => X"00000000",
		16#528c# => X"00000000",
		16#528d# => X"00000000",
		16#528e# => X"00000000",
		16#528f# => X"00000000",
		16#5290# => X"00000000",
		16#5291# => X"00000000",
		16#5292# => X"00000000",
		16#5293# => X"00000000",
		16#5294# => X"00000000",
		16#5295# => X"00000000",
		16#5296# => X"00000000",
		16#5297# => X"00000000",
		16#5298# => X"00000000",
		16#5299# => X"00000000",
		16#529a# => X"00000000",
		16#529b# => X"00000000",
		16#529c# => X"00000000",
		16#529d# => X"00000000",
		16#529e# => X"00000000",
		16#529f# => X"00000000",
		16#52a0# => X"00000000",
		16#52a1# => X"00000000",
		16#52a2# => X"00000000",
		16#52a3# => X"00000000",
		16#52a4# => X"00000000",
		16#52a5# => X"00000000",
		16#52a6# => X"00000000",
		16#52a7# => X"00000000",
		16#52a8# => X"00000000",
		16#52a9# => X"00000000",
		16#52aa# => X"00000000",
		16#52ab# => X"00000000",
		16#52ac# => X"00000000",
		16#52ad# => X"00000000",
		16#52ae# => X"00000000",
		16#52af# => X"00000000",
		16#52b0# => X"00000000",
		16#52b1# => X"00000000",
		16#52b2# => X"00000000",
		16#52b3# => X"00000000",
		16#52b4# => X"00000000",
		16#52b5# => X"00000000",
		16#52b6# => X"00000000",
		16#52b7# => X"00000000",
		16#52b8# => X"00000000",
		16#52b9# => X"00000000",
		16#52ba# => X"00000000",
		16#52bb# => X"00000000",
		16#52bc# => X"00000000",
		16#52bd# => X"00000000",
		16#52be# => X"00000000",
		16#52bf# => X"00000000",
		16#52c0# => X"00000000",
		16#52c1# => X"00000000",
		16#52c2# => X"00000000",
		16#52c3# => X"00000000",
		16#52c4# => X"00000000",
		16#52c5# => X"00000000",
		16#52c6# => X"00000000",
		16#52c7# => X"00000000",
		16#52c8# => X"00000000",
		16#52c9# => X"00000000",
		16#52ca# => X"00000000",
		16#52cb# => X"00000000",
		16#52cc# => X"00000000",
		16#52cd# => X"00000000",
		16#52ce# => X"00000000",
		16#52cf# => X"00000000",
		16#52d0# => X"00000000",
		16#52d1# => X"00000000",
		16#52d2# => X"00000000",
		16#52d3# => X"00000000",
		16#52d4# => X"00000000",
		16#52d5# => X"00000000",
		16#52d6# => X"00000000",
		16#52d7# => X"00000000",
		16#52d8# => X"00000000",
		16#52d9# => X"00000000",
		16#52da# => X"00000000",
		16#52db# => X"00000000",
		16#52dc# => X"00000000",
		16#52dd# => X"00000000",
		16#52de# => X"00000000",
		16#52df# => X"00000000",
		16#52e0# => X"00000000",
		16#52e1# => X"00000000",
		16#52e2# => X"00000000",
		16#52e3# => X"00000000",
		16#52e4# => X"00000000",
		16#52e5# => X"00000000",
		16#52e6# => X"00000000",
		16#52e7# => X"00000000",
		16#52e8# => X"00000000",
		16#52e9# => X"00000000",
		16#52ea# => X"00000000",
		16#52eb# => X"00000000",
		16#52ec# => X"00000000",
		16#52ed# => X"00000000",
		16#52ee# => X"00000000",
		16#52ef# => X"00000000",
		16#52f0# => X"00000000",
		16#52f1# => X"00000000",
		16#52f2# => X"00000000",
		16#52f3# => X"00000000",
		16#52f4# => X"00000000",
		16#52f5# => X"00000000",
		16#52f6# => X"00000000",
		16#52f7# => X"00000000",
		16#52f8# => X"00000000",
		16#52f9# => X"00000000",
		16#52fa# => X"00000000",
		16#52fb# => X"00000000",
		16#52fc# => X"00000000",
		16#52fd# => X"00000000",
		16#52fe# => X"00000000",
		16#52ff# => X"00000000",
		16#5300# => X"00000000",
		16#5301# => X"00000000",
		16#5302# => X"00000000",
		16#5303# => X"00000000",
		16#5304# => X"00000000",
		16#5305# => X"00000000",
		16#5306# => X"00000000",
		16#5307# => X"00000000",
		16#5308# => X"00000000",
		16#5309# => X"00000000",
		16#530a# => X"00000000",
		16#530b# => X"00000000",
		16#530c# => X"00000000",
		16#530d# => X"00000000",
		16#530e# => X"00000000",
		16#530f# => X"00000000",
		16#5310# => X"00000000",
		16#5311# => X"00000000",
		16#5312# => X"00000000",
		16#5313# => X"00000000",
		16#5314# => X"00000000",
		16#5315# => X"00000000",
		16#5316# => X"00000000",
		16#5317# => X"00000000",
		16#5318# => X"00000000",
		16#5319# => X"00000000",
		16#531a# => X"00000000",
		16#531b# => X"00000000",
		16#531c# => X"00000000",
		16#531d# => X"00000000",
		16#531e# => X"00000000",
		16#531f# => X"00000000",
		16#5320# => X"00000000",
		16#5321# => X"00000000",
		16#5322# => X"00000000",
		16#5323# => X"00000000",
		16#5324# => X"00000000",
		16#5325# => X"00000000",
		16#5326# => X"00000000",
		16#5327# => X"00000000",
		16#5328# => X"43000000",
		16#5329# => X"00000000",
		16#532a# => X"00000000",
		16#532b# => X"00000000",
		16#532c# => X"00000000",
		16#532d# => X"00000000",
		16#532e# => X"00000000",
		16#532f# => X"00000000",
		16#5330# => X"43000000",
		16#5331# => X"00000000",
		16#5332# => X"00000000",
		16#5333# => X"00000000",
		16#5334# => X"00000000",
		16#5335# => X"00000000",
		16#5336# => X"00000000",
		16#5337# => X"00000000",
		16#5338# => X"43000000",
		16#5339# => X"00000000",
		16#533a# => X"00000000",
		16#533b# => X"00000000",
		16#533c# => X"00000000",
		16#533d# => X"00000000",
		16#533e# => X"00000000",
		16#533f# => X"00000000",
		16#5340# => X"43000000",
		16#5341# => X"00000000",
		16#5342# => X"00000000",
		16#5343# => X"00000000",
		16#5344# => X"00000000",
		16#5345# => X"00000000",
		16#5346# => X"00000000",
		16#5347# => X"00000000",
		16#5348# => X"43000000",
		16#5349# => X"00000000",
		16#534a# => X"00000000",
		16#534b# => X"00000000",
		16#534c# => X"00000000",
		16#534d# => X"00000000",
		16#534e# => X"00000000",
		16#534f# => X"00000000",
		16#5350# => X"43000000",
		16#5351# => X"00000000",
		16#5352# => X"00000000",
		16#5353# => X"00000000",
		16#5354# => X"00000000",
		16#5355# => X"00000000",
		16#5356# => X"00000000",
		16#5357# => X"00000000",
		16#5358# => X"43000000",
		16#5359# => X"00000000",
		16#535a# => X"00000000",
		16#535b# => X"00000000",
		16#535c# => X"00000000",
		16#535d# => X"00000000",
		16#535e# => X"00000000",
		16#535f# => X"00000000",
		16#5360# => X"b4bb0010",
		16#5361# => X"20730010",
		16#5362# => X"00000000",
		16#5363# => X"78430110",
		16#5364# => X"64390110",
		16#5365# => X"743a0110",
		16#5366# => X"743a0110",
		16#5367# => X"743a0110",
		16#5368# => X"743a0110",
		16#5369# => X"743a0110",
		16#536a# => X"743a0110",
		16#536b# => X"743a0110",
		16#536c# => X"743a0110",
		16#536d# => X"743a0110",
		16#536e# => X"ffffffff",
		16#536f# => X"ffffffff",
		16#5370# => X"ffffffff",
		16#5371# => X"ffff0000",
		16#5372# => X"01004153",
		16#5373# => X"43494900",
		16#5374# => X"00000000",
		16#5375# => X"00000000",
		16#5376# => X"00000000",
		16#5377# => X"00000000",
		16#5378# => X"00000000",
		16#5379# => X"00000000",
		16#537a# => X"00004153",
		16#537b# => X"43494900",
		16#537c# => X"00000000",
		16#537d# => X"00000000",
		16#537e# => X"00000000",
		16#537f# => X"00000000",
		16#5380# => X"00000000",
		16#5381# => X"00000000",
		16#5382# => X"00000000",
		16#5383# => X"00000000",
		16#5384# => X"00000000",
		16#5385# => X"0c4e0110",
		16#5386# => X"0c4e0110",
		16#5387# => X"144e0110",
		16#5388# => X"144e0110",
		16#5389# => X"1c4e0110",
		16#538a# => X"1c4e0110",
		16#538b# => X"244e0110",
		16#538c# => X"244e0110",
		16#538d# => X"2c4e0110",
		16#538e# => X"2c4e0110",
		16#538f# => X"344e0110",
		16#5390# => X"344e0110",
		16#5391# => X"3c4e0110",
		16#5392# => X"3c4e0110",
		16#5393# => X"444e0110",
		16#5394# => X"444e0110",
		16#5395# => X"4c4e0110",
		16#5396# => X"4c4e0110",
		16#5397# => X"544e0110",
		16#5398# => X"544e0110",
		16#5399# => X"5c4e0110",
		16#539a# => X"5c4e0110",
		16#539b# => X"644e0110",
		16#539c# => X"644e0110",
		16#539d# => X"6c4e0110",
		16#539e# => X"6c4e0110",
		16#539f# => X"744e0110",
		16#53a0# => X"744e0110",
		16#53a1# => X"7c4e0110",
		16#53a2# => X"7c4e0110",
		16#53a3# => X"844e0110",
		16#53a4# => X"844e0110",
		16#53a5# => X"8c4e0110",
		16#53a6# => X"8c4e0110",
		16#53a7# => X"944e0110",
		16#53a8# => X"944e0110",
		16#53a9# => X"9c4e0110",
		16#53aa# => X"9c4e0110",
		16#53ab# => X"a44e0110",
		16#53ac# => X"a44e0110",
		16#53ad# => X"ac4e0110",
		16#53ae# => X"ac4e0110",
		16#53af# => X"b44e0110",
		16#53b0# => X"b44e0110",
		16#53b1# => X"bc4e0110",
		16#53b2# => X"bc4e0110",
		16#53b3# => X"c44e0110",
		16#53b4# => X"c44e0110",
		16#53b5# => X"cc4e0110",
		16#53b6# => X"cc4e0110",
		16#53b7# => X"d44e0110",
		16#53b8# => X"d44e0110",
		16#53b9# => X"dc4e0110",
		16#53ba# => X"dc4e0110",
		16#53bb# => X"e44e0110",
		16#53bc# => X"e44e0110",
		16#53bd# => X"ec4e0110",
		16#53be# => X"ec4e0110",
		16#53bf# => X"f44e0110",
		16#53c0# => X"f44e0110",
		16#53c1# => X"fc4e0110",
		16#53c2# => X"fc4e0110",
		16#53c3# => X"044f0110",
		16#53c4# => X"044f0110",
		16#53c5# => X"0c4f0110",
		16#53c6# => X"0c4f0110",
		16#53c7# => X"144f0110",
		16#53c8# => X"144f0110",
		16#53c9# => X"1c4f0110",
		16#53ca# => X"1c4f0110",
		16#53cb# => X"244f0110",
		16#53cc# => X"244f0110",
		16#53cd# => X"2c4f0110",
		16#53ce# => X"2c4f0110",
		16#53cf# => X"344f0110",
		16#53d0# => X"344f0110",
		16#53d1# => X"3c4f0110",
		16#53d2# => X"3c4f0110",
		16#53d3# => X"444f0110",
		16#53d4# => X"444f0110",
		16#53d5# => X"4c4f0110",
		16#53d6# => X"4c4f0110",
		16#53d7# => X"544f0110",
		16#53d8# => X"544f0110",
		16#53d9# => X"5c4f0110",
		16#53da# => X"5c4f0110",
		16#53db# => X"644f0110",
		16#53dc# => X"644f0110",
		16#53dd# => X"6c4f0110",
		16#53de# => X"6c4f0110",
		16#53df# => X"744f0110",
		16#53e0# => X"744f0110",
		16#53e1# => X"7c4f0110",
		16#53e2# => X"7c4f0110",
		16#53e3# => X"844f0110",
		16#53e4# => X"844f0110",
		16#53e5# => X"8c4f0110",
		16#53e6# => X"8c4f0110",
		16#53e7# => X"944f0110",
		16#53e8# => X"944f0110",
		16#53e9# => X"9c4f0110",
		16#53ea# => X"9c4f0110",
		16#53eb# => X"a44f0110",
		16#53ec# => X"a44f0110",
		16#53ed# => X"ac4f0110",
		16#53ee# => X"ac4f0110",
		16#53ef# => X"b44f0110",
		16#53f0# => X"b44f0110",
		16#53f1# => X"bc4f0110",
		16#53f2# => X"bc4f0110",
		16#53f3# => X"c44f0110",
		16#53f4# => X"c44f0110",
		16#53f5# => X"cc4f0110",
		16#53f6# => X"cc4f0110",
		16#53f7# => X"d44f0110",
		16#53f8# => X"d44f0110",
		16#53f9# => X"dc4f0110",
		16#53fa# => X"dc4f0110",
		16#53fb# => X"e44f0110",
		16#53fc# => X"e44f0110",
		16#53fd# => X"ec4f0110",
		16#53fe# => X"ec4f0110",
		16#53ff# => X"f44f0110",
		16#5400# => X"f44f0110",
		16#5401# => X"fc4f0110",
		16#5402# => X"fc4f0110",
		16#5403# => X"04500110",
		16#5404# => X"04500110",
		16#5405# => X"0c500110",
		16#5406# => X"0c500110",
		16#5407# => X"14500110",
		16#5408# => X"14500110",
		16#5409# => X"1c500110",
		16#540a# => X"1c500110",
		16#540b# => X"24500110",
		16#540c# => X"24500110",
		16#540d# => X"2c500110",
		16#540e# => X"2c500110",
		16#540f# => X"34500110",
		16#5410# => X"34500110",
		16#5411# => X"3c500110",
		16#5412# => X"3c500110",
		16#5413# => X"44500110",
		16#5414# => X"44500110",
		16#5415# => X"4c500110",
		16#5416# => X"4c500110",
		16#5417# => X"54500110",
		16#5418# => X"54500110",
		16#5419# => X"5c500110",
		16#541a# => X"5c500110",
		16#541b# => X"64500110",
		16#541c# => X"64500110",
		16#541d# => X"6c500110",
		16#541e# => X"6c500110",
		16#541f# => X"74500110",
		16#5420# => X"74500110",
		16#5421# => X"7c500110",
		16#5422# => X"7c500110",
		16#5423# => X"84500110",
		16#5424# => X"84500110",
		16#5425# => X"8c500110",
		16#5426# => X"8c500110",
		16#5427# => X"94500110",
		16#5428# => X"94500110",
		16#5429# => X"9c500110",
		16#542a# => X"9c500110",
		16#542b# => X"a4500110",
		16#542c# => X"a4500110",
		16#542d# => X"ac500110",
		16#542e# => X"ac500110",
		16#542f# => X"b4500110",
		16#5430# => X"b4500110",
		16#5431# => X"bc500110",
		16#5432# => X"bc500110",
		16#5433# => X"c4500110",
		16#5434# => X"c4500110",
		16#5435# => X"cc500110",
		16#5436# => X"cc500110",
		16#5437# => X"d4500110",
		16#5438# => X"d4500110",
		16#5439# => X"dc500110",
		16#543a# => X"dc500110",
		16#543b# => X"e4500110",
		16#543c# => X"e4500110",
		16#543d# => X"ec500110",
		16#543e# => X"ec500110",
		16#543f# => X"f4500110",
		16#5440# => X"f4500110",
		16#5441# => X"fc500110",
		16#5442# => X"fc500110",
		16#5443# => X"04510110",
		16#5444# => X"04510110",
		16#5445# => X"0c510110",
		16#5446# => X"0c510110",
		16#5447# => X"14510110",
		16#5448# => X"14510110",
		16#5449# => X"1c510110",
		16#544a# => X"1c510110",
		16#544b# => X"24510110",
		16#544c# => X"24510110",
		16#544d# => X"2c510110",
		16#544e# => X"2c510110",
		16#544f# => X"34510110",
		16#5450# => X"34510110",
		16#5451# => X"3c510110",
		16#5452# => X"3c510110",
		16#5453# => X"44510110",
		16#5454# => X"44510110",
		16#5455# => X"4c510110",
		16#5456# => X"4c510110",
		16#5457# => X"54510110",
		16#5458# => X"54510110",
		16#5459# => X"5c510110",
		16#545a# => X"5c510110",
		16#545b# => X"64510110",
		16#545c# => X"64510110",
		16#545d# => X"6c510110",
		16#545e# => X"6c510110",
		16#545f# => X"74510110",
		16#5460# => X"74510110",
		16#5461# => X"7c510110",
		16#5462# => X"7c510110",
		16#5463# => X"84510110",
		16#5464# => X"84510110",
		16#5465# => X"8c510110",
		16#5466# => X"8c510110",
		16#5467# => X"94510110",
		16#5468# => X"94510110",
		16#5469# => X"9c510110",
		16#546a# => X"9c510110",
		16#546b# => X"a4510110",
		16#546c# => X"a4510110",
		16#546d# => X"ac510110",
		16#546e# => X"ac510110",
		16#546f# => X"b4510110",
		16#5470# => X"b4510110",
		16#5471# => X"bc510110",
		16#5472# => X"bc510110",
		16#5473# => X"c4510110",
		16#5474# => X"c4510110",
		16#5475# => X"cc510110",
		16#5476# => X"cc510110",
		16#5477# => X"d4510110",
		16#5478# => X"d4510110",
		16#5479# => X"dc510110",
		16#547a# => X"dc510110",
		16#547b# => X"e4510110",
		16#547c# => X"e4510110",
		16#547d# => X"ec510110",
		16#547e# => X"ec510110",
		16#547f# => X"f4510110",
		16#5480# => X"f4510110",
		16#5481# => X"fc510110",
		16#5482# => X"fc510110",
		16#5483# => X"04520110",
		16#5484# => X"04520110",
		16#5485# => X"00000000",
		16#5486# => X"00000000",
		16#5487# => X"0000f03f",
		16#5488# => X"00000000",
		16#5489# => X"00002440",
		16#548a# => X"00000000",
		16#548b# => X"00005043",
		16#548c# => X"78480110",
		16#548d# => X"78480110",
		16#548e# => X"ffffffff",
		16#548f# => X"00000200",
		16#5490# => X"64520110",
		16#5491# => X"05000090",
		16#5492# => X"00000090",
		16#5493# => X"00000000",
		16#5494# => X"00000000",
		16#5495# => X"00000000",
		16#5496# => X"00000000",
		16#5497# => X"00000000",
		16#5498# => X"00000000",
		16#5499# => X"00000000",
		16#549a# => X"00000000",
		16#549b# => X"00000000",
		16#549c# => X"00000000",
		16#549d# => X"00000000",
		16#549e# => X"00000000",
		16#549f# => X"00000000",
		16#54a0# => X"00000000",
		16#54a1# => X"00000000",
		16#54a2# => X"00000000",
		16#54a3# => X"00000000",
		16#54a4# => X"00000000",
		16#54a5# => X"00000000",
		16#54a6# => X"00000000",
		16#54a7# => X"00000000",
		16#54a8# => X"00000000",
		16#54a9# => X"00000000",
		16#54aa# => X"00000000",
		16#54ab# => X"00000000",
		16#54ac# => X"00000000",
		16#54ad# => X"00000000",
		16#54ae# => X"00000000",
		16#54af# => X"00000000",
		16#54b0# => X"00000000",
		16#54b1# => X"00000000",
		16#54b2# => X"00000000",
		16#54b3# => X"00000000",
		16#54b4# => X"00000000",
		16#54b5# => X"00000000",
		16#54b6# => X"00000000",
		16#54b7# => X"00000000",
		16#54b8# => X"00000000",
		16#54b9# => X"00000000",
		16#54ba# => X"00000000",
		16#54bb# => X"00000000",
		16#54bc# => X"00000000",
		16#54bd# => X"00000000",
		16#54be# => X"00000000",
		16#54bf# => X"00000000",
		16#54c0# => X"00000000",
		16#54c1# => X"00000000",
		16#54c2# => X"00000000",
		16#54c3# => X"00000000",
		16#54c4# => X"00000000",
		16#54c5# => X"00000000",
		16#54c6# => X"00000000",
		16#54c7# => X"00000000",
		16#54c8# => X"00000000",
		16#54c9# => X"00000000",
		16#54ca# => X"00000000",
		16#54cb# => X"00000000",
		16#54cc# => X"00000000",
		16#54cd# => X"00000000",
		16#54ce# => X"00000000",
		16#54cf# => X"00000000",
		16#54d0# => X"00000000",
		16#54d1# => X"00000000",
		16#54d2# => X"00000000",
		16#54d3# => X"00000000",
		16#54d4# => X"00000000",
		16#54d5# => X"00000000",
		16#54d6# => X"00000000",
		16#54d7# => X"00000000",
		16#54d8# => X"00000000",
		16#54d9# => X"00000000",
		16#54da# => X"00000000",
		16#54db# => X"00000000",
		16#54dc# => X"00000000",
		16#54dd# => X"00000000",
		16#54de# => X"00000000",
		16#54df# => X"00000000",
		16#54e0# => X"00000000",
		16#54e1# => X"00000000",
		16#54e2# => X"00000000",
		16#54e3# => X"00000000",
		16#54e4# => X"00000000",
		16#54e5# => X"00000000",
		16#54e6# => X"00000000",
		16#54e7# => X"00000000",
		16#54e8# => X"00000000",
		16#54e9# => X"00000000",
		16#54ea# => X"00000000",
		16#54eb# => X"00000000",
		16#54ec# => X"00000000",
		16#54ed# => X"00000000",
		16#54ee# => X"00000000",
		16#54ef# => X"00000000",
		16#54f0# => X"00000000",
		16#54f1# => X"00000000",
		16#54f2# => X"00000000",
		16#54f3# => X"00000000",
		16#54f4# => X"00000000",
		16#54f5# => X"00000000",
		16#54f6# => X"00000000",
		16#54f7# => X"00000000",
		16#54f8# => X"00000000",
		16#54f9# => X"00000000",
		16#54fa# => X"00000000",
		16#54fb# => X"00000000",
		16#54fc# => X"00000000",
		16#54fd# => X"00000000",
		16#54fe# => X"00000000",
		16#54ff# => X"00000000",
		16#5500# => X"00000000",
		16#5501# => X"00000000",
		16#5502# => X"00000000",
		16#5503# => X"00000000",
		16#5504# => X"00000000",
		16#5505# => X"00000000",
		16#5506# => X"00000000",
		16#5507# => X"00000000",
		16#5508# => X"00000000",
		16#5509# => X"00000000",
		16#550a# => X"00000000",
		16#550b# => X"00000000",
		16#550c# => X"00000000",
		16#550d# => X"00000000",
		16#550e# => X"00000000",
		16#550f# => X"00000000",
		16#5510# => X"00000000",
		16#5511# => X"00000000",
		16#5512# => X"00000000",
		16#5513# => X"00000000",
		16#5514# => X"00000000",
		16#5515# => X"00000000",
		16#5516# => X"00000000",
		16#5517# => X"00000000",
		16#5518# => X"00000000",
		16#5519# => X"00000000",
		16#551a# => X"00000000",
		16#551b# => X"00000000",
		16#551c# => X"00000000",
		16#551d# => X"00000000",
		16#551e# => X"00000000",
		16#551f# => X"00000000",
		16#5520# => X"00000000",
		16#5521# => X"00000000",
		16#5522# => X"00000000",
		16#5523# => X"00000000",
		16#5524# => X"00000000",
		16#5525# => X"00000000",
		16#5526# => X"00000000",
		16#5527# => X"00000000",
		16#5528# => X"00000000",
		16#5529# => X"00000000",
		16#552a# => X"00000000",
		16#552b# => X"00000000",
		16#552c# => X"00000000",
		16#552d# => X"00000000",
		16#552e# => X"00000000",
		16#552f# => X"00000000",
		16#5530# => X"00000000",
		16#5531# => X"00000000",
		16#5532# => X"00000000",
		16#5533# => X"00000000",
		16#5534# => X"00000000",
		16#5535# => X"00000000",
		16#5536# => X"00000000",
		16#5537# => X"00000000",
		16#5538# => X"00000000",
		16#5539# => X"00000000",
		16#553a# => X"00000000",
		16#553b# => X"00000000",
		16#553c# => X"00000000",
		16#553d# => X"00000000",
		16#553e# => X"00000000",
		16#553f# => X"00000000",
		16#5540# => X"00000000",
		16#5541# => X"00000000",
		16#5542# => X"00000000",
		16#5543# => X"00000000",
		16#5544# => X"00000000",
		16#5545# => X"00000000",
		16#5546# => X"00000000",
		16#5547# => X"00000000",
		16#5548# => X"00000000",
		16#5549# => X"00000000",
		16#554a# => X"00000000",
		16#554b# => X"00000000",
		16#554c# => X"00000000",
		16#554d# => X"00000000",
		16#554e# => X"00000000",
		16#554f# => X"00000000",
		16#5550# => X"00000000",
		16#5551# => X"00000000",
		16#5552# => X"00000000",
		16#5553# => X"00000000",
		16#5554# => X"00000000",
		16#5555# => X"00000000",
		16#5556# => X"00000000",
		16#5557# => X"00000000",
		16#5558# => X"00000000",
		16#5559# => X"00000000",
		16#555a# => X"00000000",
		16#555b# => X"00000000",
		16#555c# => X"00000000",
		16#555d# => X"00000000",
		16#555e# => X"00000000",
		16#555f# => X"00000000",
		16#5560# => X"00000000",
		16#5561# => X"00000000",
		16#5562# => X"00000000",
		16#5563# => X"00000000",
		16#5564# => X"00000000",
		16#5565# => X"00000000",
		16#5566# => X"00000000",
		16#5567# => X"00000000",
		16#5568# => X"00000000",
		16#5569# => X"00000000",
		16#556a# => X"00000000",
		16#556b# => X"00000000",
		16#556c# => X"00000000",
		16#556d# => X"00000000",
		16#556e# => X"00000000",
		16#556f# => X"00000000",
		16#5570# => X"00000000",
		16#5571# => X"00000000",
		16#5572# => X"00000000",
		16#5573# => X"00000000",
		16#5574# => X"00000000",
		16#5575# => X"00000000",
		16#5576# => X"00000000",
		16#5577# => X"00000000",
		16#5578# => X"00000000",
		16#5579# => X"00000000",
		16#557a# => X"00000000",
		16#557b# => X"00000000",
		16#557c# => X"00000000",
		16#557d# => X"00000000",
		16#557e# => X"00000000",
		16#557f# => X"00000000",
		16#5580# => X"00000000",
		16#5581# => X"00000000",
		16#5582# => X"00000000",
		16#5583# => X"00000000",
		16#5584# => X"00000000",
		16#5585# => X"00000000",
		16#5586# => X"00000000",
		16#5587# => X"00000000",
		16#5588# => X"00000000",
		16#5589# => X"00000000",
		16#558a# => X"00000000",
		16#558b# => X"00000000",
		16#558c# => X"00000000",
		16#558d# => X"00000000",
		16#558e# => X"00000000",
		16#558f# => X"00000000",
		16#5590# => X"00000000",
		16#5591# => X"00000000",
		16#5592# => X"00000000",
		16#5593# => X"00000000",
		16#5594# => X"00000000",
		16#5595# => X"00000000",
		16#5596# => X"00000000",
		16#5597# => X"00000000",
		16#5598# => X"00000000",
		16#5599# => X"00000000",
		16#559a# => X"00000000",
		16#559b# => X"00000000",
		16#559c# => X"00000000",
		16#559d# => X"00000000",
		16#559e# => X"00000000",
		16#559f# => X"00000000",
		16#55a0# => X"00000000",
		16#55a1# => X"00000000",
		16#55a2# => X"00000000",
		16#55a3# => X"00000000",
		16#55a4# => X"00000000",
		16#55a5# => X"00000000",
		16#55a6# => X"00000000",
		16#55a7# => X"00000000",
		16#55a8# => X"00000000",
		16#55a9# => X"00000000",
		16#55aa# => X"00000000",
		16#55ab# => X"00000000",
		16#55ac# => X"00000000",
		16#55ad# => X"00000000",
		16#55ae# => X"00000000",
		16#55af# => X"00000000",
		16#55b0# => X"00000000",
		16#55b1# => X"00000000",
		16#55b2# => X"00000000",
		16#55b3# => X"00000000",
		16#55b4# => X"00000000",
		16#55b5# => X"00000000",
		16#55b6# => X"00000000",
		16#55b7# => X"00000000",
		16#55b8# => X"00000000",
		16#55b9# => X"00000000",
		16#55ba# => X"00000000",
		16#55bb# => X"00000000",
		16#55bc# => X"00000000",
		16#55bd# => X"00000000",
		16#55be# => X"00000000",
		16#55bf# => X"00000000",
		16#55c0# => X"00000000",
		16#55c1# => X"00000000",
		16#55c2# => X"00000000",
		16#55c3# => X"00000000",
		16#55c4# => X"00000000",
		16#55c5# => X"00000000",
		16#55c6# => X"00000000",
		16#55c7# => X"00000000",
		16#55c8# => X"00000000",
		16#55c9# => X"00000000",
		16#55ca# => X"00000000",
		16#55cb# => X"00000000",
		16#55cc# => X"00000000",
		16#55cd# => X"00000000",
		16#55ce# => X"00000000",
		16#55cf# => X"00000000",
		16#55d0# => X"00000000",
		16#55d1# => X"00000000",
		16#55d2# => X"00000000",
		16#55d3# => X"00000000",
		16#55d4# => X"00000000",
		16#55d5# => X"00000000",
		16#55d6# => X"00000000",
		16#55d7# => X"00000000",
		16#55d8# => X"00000000",
		16#55d9# => X"00000000",
		16#55da# => X"00000000",
		16#55db# => X"00000000",
		16#55dc# => X"00000000",
		16#55dd# => X"00000000",
		16#55de# => X"00000000",
		16#55df# => X"00000000",
		16#55e0# => X"00000000",
		16#55e1# => X"00000000",
		16#55e2# => X"00000000",
		16#55e3# => X"00000000",
		16#55e4# => X"00000000",
		16#55e5# => X"00000000",
		16#55e6# => X"00000000",
		16#55e7# => X"00000000",
		16#55e8# => X"00000000",
		16#55e9# => X"00000000",
		16#55ea# => X"00000000",
		16#55eb# => X"00000000",
		16#55ec# => X"00000000",
		16#55ed# => X"00000000",
		16#55ee# => X"00000000",
		16#55ef# => X"00000000",
		16#55f0# => X"00000000",
		16#55f1# => X"00000000",
		16#55f2# => X"00000000",
		16#55f3# => X"00000000",
		16#55f4# => X"00000000",
		16#55f5# => X"00000000",
		16#55f6# => X"00000000",
		16#55f7# => X"00000000",
		16#55f8# => X"00000000",
		16#55f9# => X"00000000",
		16#55fa# => X"00000000",
		16#55fb# => X"00000000",
		16#55fc# => X"00000000",
		16#55fd# => X"00000000",
		16#55fe# => X"00000000",
		16#55ff# => X"00000000",
		16#5600# => X"00000000",
		16#5601# => X"00000000",
		16#5602# => X"00000000",
		16#5603# => X"00000000",
		16#5604# => X"00000000",
		16#5605# => X"00000000",
		16#5606# => X"00000000",
		16#5607# => X"00000000",
		16#5608# => X"00000000",
		16#5609# => X"00000000",
		16#560a# => X"00000000",
		16#560b# => X"00000000",
		16#560c# => X"00000000",
		16#560d# => X"00000000",
		16#560e# => X"00000000",
		16#560f# => X"00000000",
		16#5610# => X"00000000",
		16#5611# => X"00000000",
		16#5612# => X"00000000",
		16#5613# => X"00000000",
		16#5614# => X"00000000",
		16#5615# => X"00000000",
		16#5616# => X"00000000",
		16#5617# => X"00000000",
		16#5618# => X"00000000",
		16#5619# => X"00000000",
		16#561a# => X"00000000",
		16#561b# => X"00000000",
		16#561c# => X"00000000",
		16#561d# => X"00000000",
		16#561e# => X"00000000",
		16#561f# => X"00000000",
		16#5620# => X"00000000",
		16#5621# => X"00000000",
		16#5622# => X"00000000",
		16#5623# => X"00000000",
		16#5624# => X"00000000",
		16#5625# => X"00000000",
		16#5626# => X"00000000",
		16#5627# => X"00000000",
		16#5628# => X"00000000",
		16#5629# => X"00000000",
		16#562a# => X"00000000",
		16#562b# => X"00000000",
		16#562c# => X"00000000",
		16#562d# => X"00000000",
		16#562e# => X"00000000",
		16#562f# => X"00000000",
		16#5630# => X"00000000",
		16#5631# => X"00000000",
		16#5632# => X"00000000",
		16#5633# => X"00000000",
		16#5634# => X"00000000",
		16#5635# => X"00000000",
		16#5636# => X"00000000",
		16#5637# => X"00000000",
		16#5638# => X"00000000",
		16#5639# => X"00000000",
		16#563a# => X"00000000",
		16#563b# => X"00000000",
		16#563c# => X"00000000",
		16#563d# => X"00000000",
		16#563e# => X"00000000",
		16#563f# => X"00000000",
		16#5640# => X"00000000",
		16#5641# => X"00000000",
		16#5642# => X"00000000",
		16#5643# => X"00000000",
		16#5644# => X"00000000",
		16#5645# => X"00000000",
		16#5646# => X"00000000",
		16#5647# => X"00000000",
		16#5648# => X"00000000",
		16#5649# => X"00000000",
		16#564a# => X"00000000",
		16#564b# => X"00000000",
		16#564c# => X"00000000",
		16#564d# => X"00000000",
		16#564e# => X"00000000",
		16#564f# => X"00000000",
		16#5650# => X"00000000",
		16#5651# => X"00000000",
		16#5652# => X"00000000",
		16#5653# => X"00000000",
		16#5654# => X"00000000",
		16#5655# => X"00000000",
		16#5656# => X"00000000",
		16#5657# => X"00000000",
		16#5658# => X"00000000",
		16#5659# => X"00000000",
		16#565a# => X"00000000",
		16#565b# => X"00000000",
		16#565c# => X"00000000",
		16#565d# => X"00000000",
		16#565e# => X"00000000",
		16#565f# => X"00000000",
		16#5660# => X"00000000",
		16#5661# => X"00000000",
		16#5662# => X"00000000",
		16#5663# => X"00000000",
		16#5664# => X"00000000",
		16#5665# => X"00000000",
		16#5666# => X"00000000",
		16#5667# => X"00000000",
		16#5668# => X"00000000",
		16#5669# => X"00000000",
		16#566a# => X"00000000",
		16#566b# => X"00000000",
		16#566c# => X"00000000",
		16#566d# => X"00000000",
		16#566e# => X"00000000",
		16#566f# => X"00000000",
		16#5670# => X"00000000",
		16#5671# => X"00000000",
		16#5672# => X"00000000",
		16#5673# => X"00000000",
		16#5674# => X"00000000",
		16#5675# => X"00000000",
		16#5676# => X"00000000",
		16#5677# => X"00000000",
		16#5678# => X"00000000",
		16#5679# => X"00000000",
		16#567a# => X"00000000",
		16#567b# => X"00000000",
		16#567c# => X"00000000",
		16#567d# => X"00000000",
		16#567e# => X"00000000",
		16#567f# => X"00000000",
		16#5680# => X"00000000",
		16#5681# => X"00000000",
		16#5682# => X"00000000",
		16#5683# => X"00000000",
		16#5684# => X"00000000",
		16#5685# => X"00000000",
		16#5686# => X"00000000",
		16#5687# => X"00000000",
		16#5688# => X"00000000",
		16#5689# => X"00000000",
		16#568a# => X"00000000",
		16#568b# => X"00000000",
		16#568c# => X"00000000",
		16#568d# => X"00000000",
		16#568e# => X"00000000",
		16#568f# => X"00000000",
		16#5690# => X"00000000",
		16#5691# => X"00000000",
		16#5692# => X"00000000",
		16#5693# => X"00000000",
		16#5694# => X"00000000",
		16#5695# => X"00000000",
		16#5696# => X"00000000",
		16#5697# => X"00000000",
		16#5698# => X"00000000",
		16#5699# => X"00000000",
		16#569a# => X"00000000",
		16#569b# => X"00000000",
		16#569c# => X"00000000",
		16#569d# => X"00000000",
		16#569e# => X"00000000",
		16#569f# => X"00000000",
		16#56a0# => X"00000000",
		16#56a1# => X"00000000",
		16#56a2# => X"00000000",
		16#56a3# => X"00000000",
		16#56a4# => X"00000000",
		16#56a5# => X"00000000",
		16#56a6# => X"00000000",
		16#56a7# => X"00000000",
		16#56a8# => X"00000000",
		16#56a9# => X"00000000",
		16#56aa# => X"00000000",
		16#56ab# => X"00000000",
		16#56ac# => X"00000000",
		16#56ad# => X"00000000",
		16#56ae# => X"00000000",
		16#56af# => X"00000000",
		16#56b0# => X"00000000",
		16#56b1# => X"00000000",
		16#56b2# => X"00000000",
		16#56b3# => X"00000000",
		16#56b4# => X"00000000",
		16#56b5# => X"00000000",
		16#56b6# => X"00000000",
		16#56b7# => X"00000000",
		16#56b8# => X"00000000",
		16#56b9# => X"00000000",
		16#56ba# => X"00000000",
		16#56bb# => X"00000000",
		16#56bc# => X"00000000",
		16#56bd# => X"00000000",
		16#56be# => X"00000000",
		16#56bf# => X"00000000",
		16#56c0# => X"00000000",
		16#56c1# => X"00000000",
		16#56c2# => X"00000000",
		16#56c3# => X"00000000",
		16#56c4# => X"00000000",
		16#56c5# => X"00000000",
		16#56c6# => X"00000000",
		16#56c7# => X"00000000",
		16#56c8# => X"00000000",
		16#56c9# => X"00000000",
		16#56ca# => X"00000000",
		16#56cb# => X"00000000",
		16#56cc# => X"00000000",
		16#56cd# => X"00000000",
		16#56ce# => X"00000000",
		16#56cf# => X"00000000",
		16#56d0# => X"00000000",
		16#56d1# => X"00000000",
		16#56d2# => X"00000000",
		16#56d3# => X"00000000",
		16#56d4# => X"00000000",
		16#56d5# => X"00000000",
		16#56d6# => X"00000000",
		16#56d7# => X"00000000",
		16#56d8# => X"00000000",
		16#56d9# => X"00000000",
		16#56da# => X"00000000",
		16#56db# => X"00000000",
		16#56dc# => X"00000000",
		16#56dd# => X"00000000",
		16#56de# => X"00000000",
		16#56df# => X"00000000",
		16#56e0# => X"00000000",
		16#56e1# => X"00000000",
		16#56e2# => X"00000000",
		16#56e3# => X"00000000",
		16#56e4# => X"00000000",
		16#56e5# => X"00000000",
		16#56e6# => X"00000000",
		16#56e7# => X"00000000",
		16#56e8# => X"00000000",
		16#56e9# => X"00000000",
		16#56ea# => X"00000000",
		16#56eb# => X"00000000",
		16#56ec# => X"00000000",
		16#56ed# => X"00000000",
		16#56ee# => X"00000000",
		16#56ef# => X"00000000",
		16#56f0# => X"00000000",
		16#56f1# => X"00000000",
		16#56f2# => X"00000000",
		16#56f3# => X"00000000",
		16#56f4# => X"00000000",
		16#56f5# => X"00000000",
		16#56f6# => X"00000000",
		16#56f7# => X"00000000",
		16#56f8# => X"00000000",
		16#56f9# => X"00000000",
		16#56fa# => X"00000000",
		16#56fb# => X"00000000",
		16#56fc# => X"00000000",
		16#56fd# => X"00000000",
		16#56fe# => X"00000000",
		16#56ff# => X"00000000",
		16#5700# => X"00000000",
		16#5701# => X"00000000",
		16#5702# => X"00000000",
		16#5703# => X"00000000",
		16#5704# => X"00000000",
		16#5705# => X"00000000",
		16#5706# => X"00000000",
		16#5707# => X"00000000",
		16#5708# => X"00000000",
		16#5709# => X"00000000",
		16#570a# => X"00000000",
		16#570b# => X"00000000",
		16#570c# => X"00000000",
		16#570d# => X"00000000",
		16#570e# => X"00000000",
		16#570f# => X"00000000",
		16#5710# => X"00000000",
		16#5711# => X"00000000",
		16#5712# => X"00000000",
		16#5713# => X"00000000",
		16#5714# => X"00000000",
		16#5715# => X"00000000",
		16#5716# => X"00000000",
		16#5717# => X"00000000",
		16#5718# => X"00000000",
		16#5719# => X"00000000",
		16#571a# => X"00000000",
		16#571b# => X"00000000",
		16#571c# => X"00000000",
		16#571d# => X"00000000",
		16#571e# => X"00000000",
		16#571f# => X"00000000",
		16#5720# => X"00000000",
		16#5721# => X"00000000",
		16#5722# => X"00000000",
		16#5723# => X"00000000",
		16#5724# => X"00000000",
		16#5725# => X"00000000",
		16#5726# => X"00000000",
		16#5727# => X"00000000",
		16#5728# => X"00000000",
		16#5729# => X"00000000",
		16#572a# => X"00000000",
		16#572b# => X"00000000",
		16#572c# => X"00000000",
		16#572d# => X"00000000",
		16#572e# => X"00000000",
		16#572f# => X"00000000",
		16#5730# => X"00000000",
		16#5731# => X"00000000",
		16#5732# => X"00000000",
		16#5733# => X"00000000",
		16#5734# => X"00000000",
		16#5735# => X"00000000",
		16#5736# => X"00000000",
		16#5737# => X"00000000",
		16#5738# => X"00000000",
		16#5739# => X"00000000",
		16#573a# => X"00000000",
		16#573b# => X"00000000",
		16#573c# => X"00000000",
		16#573d# => X"00000000",
		16#573e# => X"00000000",
		16#573f# => X"00000000",
		16#5740# => X"00000000",
		16#5741# => X"00000000",
		16#5742# => X"00000000",
		16#5743# => X"00000000",
		16#5744# => X"00000000",
		16#5745# => X"00000000",
		16#5746# => X"00000000",
		16#5747# => X"00000000",
		16#5748# => X"00000000",
		16#5749# => X"00000000",
		16#574a# => X"00000000",
		16#574b# => X"00000000",
		16#574c# => X"00000000",
		16#574d# => X"00000000",
		16#574e# => X"00000000",
		16#574f# => X"00000000",
		16#5750# => X"00000000",
		16#5751# => X"00000000",
		16#5752# => X"00000000",
		16#5753# => X"00000000",
		16#5754# => X"00000000",
		16#5755# => X"00000000",
		16#5756# => X"00000000",
		16#5757# => X"00000000",
		16#5758# => X"00000000",
		16#5759# => X"00000000",
		16#575a# => X"00000000",
		16#575b# => X"00000000",
		16#575c# => X"00000000",
		16#575d# => X"00000000",
		16#575e# => X"00000000",
		16#575f# => X"00000000",
		16#5760# => X"00000000",
		16#5761# => X"00000000",
		16#5762# => X"00000000",
		16#5763# => X"00000000",
		16#5764# => X"00000000",
		16#5765# => X"00000000",
		16#5766# => X"00000000",
		16#5767# => X"00000000",
		16#5768# => X"00000000",
		16#5769# => X"00000000",
		16#576a# => X"00000000",
		16#576b# => X"00000000",
		16#576c# => X"00000000",
		16#576d# => X"00000000",
		16#576e# => X"00000000",
		16#576f# => X"00000000",
		16#5770# => X"00000000",
		16#5771# => X"00000000",
		16#5772# => X"00000000",
		16#5773# => X"00000000",
		16#5774# => X"00000000",
		16#5775# => X"00000000",
		16#5776# => X"00000000",
		16#5777# => X"00000000",
		16#5778# => X"00000000",
		16#5779# => X"00000000",
		16#577a# => X"00000000",
		16#577b# => X"00000000",
		16#577c# => X"00000000",
		16#577d# => X"00000000",
		16#577e# => X"00000000",
		16#577f# => X"00000000",
		16#5780# => X"00000000",
		16#5781# => X"00000000",
		16#5782# => X"00000000",
		16#5783# => X"00000000",
		16#5784# => X"00000000",
		16#5785# => X"00000000",
		16#5786# => X"00000000",
		16#5787# => X"00000000",
		16#5788# => X"00000000",
		16#5789# => X"00000000",
		16#578a# => X"00000000",
		16#578b# => X"00000000",
		16#578c# => X"00000000",
		16#578d# => X"00000000",
		16#578e# => X"00000000",
		16#578f# => X"00000000",
		16#5790# => X"00000000",
		16#5791# => X"00000000",
		16#5792# => X"00000000",
		16#5793# => X"00000000",
		16#5794# => X"00000000",
		16#5795# => X"00000000",
		16#5796# => X"00000000",
		16#5797# => X"00000000",
		16#5798# => X"00000000",
		16#5799# => X"00000000",
		16#579a# => X"00000000",
		16#579b# => X"00000000",
		16#579c# => X"00000000",
		16#579d# => X"00000000",
		16#579e# => X"00000000",
		16#579f# => X"00000000",
		16#57a0# => X"00000000",
		16#57a1# => X"00000000",
		16#57a2# => X"00000000",
		16#57a3# => X"00000000",
		16#57a4# => X"00000000",
		16#57a5# => X"00000000",
		16#57a6# => X"00000000",
		16#57a7# => X"00000000",
		16#57a8# => X"00000000",
		16#57a9# => X"00000000",
		16#57aa# => X"00000000",
		16#57ab# => X"00000000",
		16#57ac# => X"00000000",
		16#57ad# => X"00000000",
		16#57ae# => X"00000000",
		16#57af# => X"00000000",
		16#57b0# => X"00000000",
		16#57b1# => X"00000000",
		16#57b2# => X"00000000",
		16#57b3# => X"00000000",
		16#57b4# => X"00000000",
		16#57b5# => X"00000000",
		16#57b6# => X"00000000",
		16#57b7# => X"00000000",
		16#57b8# => X"00000000",
		16#57b9# => X"00000000",
		16#57ba# => X"00000000",
		16#57bb# => X"00000000",
		16#57bc# => X"00000000",
		16#57bd# => X"00000000",
		16#57be# => X"00000000",
		16#57bf# => X"00000000",
		16#57c0# => X"00000000",
		16#57c1# => X"00000000",
		16#57c2# => X"00000000",
		16#57c3# => X"00000000",
		16#57c4# => X"00000000",
		16#57c5# => X"00000000",
		16#57c6# => X"00000000",
		16#57c7# => X"00000000",
		16#57c8# => X"00000000",
		16#57c9# => X"00000000",
		16#57ca# => X"00000000",
		16#57cb# => X"00000000",
		16#57cc# => X"00000000",
		16#57cd# => X"00000000",
		16#57ce# => X"00000000",
		16#57cf# => X"00000000",
		16#57d0# => X"00000000",
		16#57d1# => X"00000000",
		16#57d2# => X"00000000",
		16#57d3# => X"00000000",
		16#57d4# => X"00000000",
		16#57d5# => X"00000000",
		16#57d6# => X"00000000",
		16#57d7# => X"00000000",
		16#57d8# => X"00000000",
		16#57d9# => X"00000000",
		16#57da# => X"00000000",
		16#57db# => X"00000000",
		16#57dc# => X"00000000",
		16#57dd# => X"00000000",
		16#57de# => X"00000000",
		16#57df# => X"00000000",
		16#57e0# => X"00000000",
		16#57e1# => X"00000000",
		16#57e2# => X"00000000",
		16#57e3# => X"00000000",
		16#57e4# => X"00000000",
		16#57e5# => X"00000000",
		16#57e6# => X"00000000",
		16#57e7# => X"00000000",
		16#57e8# => X"00000000",
		16#57e9# => X"00000000",
		16#57ea# => X"00000000",
		16#57eb# => X"00000000",
		16#57ec# => X"00000000",
		16#57ed# => X"00000000",
		16#57ee# => X"00000000",
		16#57ef# => X"00000000",
		16#57f0# => X"00000000",
		16#57f1# => X"00000000",
		16#57f2# => X"00000000",
		16#57f3# => X"00000000",
		16#57f4# => X"00000000",
		16#57f5# => X"00000000",
		16#57f6# => X"00000000",
		16#57f7# => X"00000000",
		16#57f8# => X"00000000",
		16#57f9# => X"00000000",
		16#57fa# => X"00000000",
		16#57fb# => X"00000000",
		16#57fc# => X"00000000",
		16#57fd# => X"00000000",
		16#57fe# => X"00000000",
		16#57ff# => X"00000000",
		16#5800# => X"00000000",
		16#5801# => X"00000000",
		16#5802# => X"00000000",
		16#5803# => X"00000000",
		16#5804# => X"00000000",
		16#5805# => X"00000000",
		16#5806# => X"00000000",
		16#5807# => X"00000000",
		16#5808# => X"00000000",
		16#5809# => X"00000000",
		16#580a# => X"00000000",
		16#580b# => X"00000000",
		16#580c# => X"00000000",
		16#580d# => X"00000000",
		16#580e# => X"00000000",
		16#580f# => X"00000000",
		16#5810# => X"00000000",
		16#5811# => X"00000000",
		16#5812# => X"00000000",
		16#5813# => X"00000000",
		16#5814# => X"00000000",
		16#5815# => X"00000000",
		16#5816# => X"00000000",
		16#5817# => X"00000000",
		16#5818# => X"00000000",
		16#5819# => X"00000000",
		16#581a# => X"00000000",
		16#581b# => X"00000000",
		16#581c# => X"00000000",
		16#581d# => X"00000000",
		16#581e# => X"00000000",
		16#581f# => X"00000000",
		16#5820# => X"00000000",
		16#5821# => X"00000000",
		16#5822# => X"00000000",
		16#5823# => X"00000000",
		16#5824# => X"00000000",
		16#5825# => X"00000000",
		16#5826# => X"00000000",
		16#5827# => X"00000000",
		16#5828# => X"00000000",
		16#5829# => X"00000000",
		16#582a# => X"00000000",
		16#582b# => X"00000000",
		16#582c# => X"00000000",
		16#582d# => X"00000000",
		16#582e# => X"00000000",
		16#582f# => X"00000000",
		16#5830# => X"00000000",
		16#5831# => X"00000000",
		16#5832# => X"00000000",
		16#5833# => X"00000000",
		16#5834# => X"00000000",
		16#5835# => X"00000000",
		16#5836# => X"00000000",
		16#5837# => X"00000000",
		16#5838# => X"00000000",
		16#5839# => X"00000000",
		16#583a# => X"00000000",
		16#583b# => X"00000000",
		16#583c# => X"00000000",
		16#583d# => X"00000000",
		16#583e# => X"00000000",
		16#583f# => X"00000000",
		16#5840# => X"00000000",
		16#5841# => X"00000000",
		16#5842# => X"00000000",
		16#5843# => X"00000000",
		16#5844# => X"00000000",
		16#5845# => X"00000000",
		16#5846# => X"00000000",
		16#5847# => X"00000000",
		16#5848# => X"00000000",
		16#5849# => X"00000000",
		16#584a# => X"00000000",
		16#584b# => X"00000000",
		16#584c# => X"00000000",
		16#584d# => X"00000000",
		16#584e# => X"00000000",
		16#584f# => X"00000000",
		16#5850# => X"00000000",
		16#5851# => X"00000000",
		16#5852# => X"00000000",
		16#5853# => X"00000000",
		16#5854# => X"00000000",
		16#5855# => X"00000000",
		16#5856# => X"00000000",
		16#5857# => X"00000000",
		16#5858# => X"00000000",
		16#5859# => X"00000000",
		16#585a# => X"00000000",
		16#585b# => X"00000000",
		16#585c# => X"00000000",
		16#585d# => X"00000000",
		16#585e# => X"00000000",
		16#585f# => X"00000000",
		16#5860# => X"00000000",
		16#5861# => X"00000000",
		16#5862# => X"00000000",
		16#5863# => X"00000000",
		16#5864# => X"00000000",
		16#5865# => X"00000000",
		16#5866# => X"00000000",
		16#5867# => X"00000000",
		16#5868# => X"00000000",
		16#5869# => X"00000000",
		16#586a# => X"00000000",
		16#586b# => X"00000000",
		16#586c# => X"00000000",
		16#586d# => X"00000000",
		16#586e# => X"00000000",
		16#586f# => X"00000000",
		16#5870# => X"00000000",
		16#5871# => X"00000000",
		16#5872# => X"00000000",
		16#5873# => X"00000000",
		16#5874# => X"00000000",
		16#5875# => X"00000000",
		16#5876# => X"00000000",
		16#5877# => X"00000000",
		16#5878# => X"00000000",
		16#5879# => X"00000000",
		16#587a# => X"00000000",
		16#587b# => X"00000000",
		16#587c# => X"00000000",
		16#587d# => X"00000000",
		16#587e# => X"00000000",
		16#587f# => X"00000000",
		16#5880# => X"00000000",
		16#5881# => X"00000000",
		16#5882# => X"00000000",
		16#5883# => X"00000000",
		16#5884# => X"00000000",
		16#5885# => X"00000000",
		16#5886# => X"00000000",
		16#5887# => X"00000000",
		16#5888# => X"00000000",
		16#5889# => X"00000000",
		16#588a# => X"00000000",
		16#588b# => X"00000000",
		16#588c# => X"00000000",
		16#588d# => X"00000000",
		16#588e# => X"00000000",
		16#588f# => X"00000000",
		16#5890# => X"00000000",
		16#5891# => X"00000000",
		16#5892# => X"00000000",
		16#5893# => X"00000000",
		16#5894# => X"00000000",
		16#5895# => X"00000000",
		16#5896# => X"00000000",
		16#5897# => X"00000000",
		16#5898# => X"00000000",
		16#5899# => X"00000000",
		16#589a# => X"00000000",
		16#589b# => X"00000000",
		16#589c# => X"00000000",
		16#589d# => X"00000000",
		16#589e# => X"00000000",
		16#589f# => X"00000000",
		16#58a0# => X"00000000",
		16#58a1# => X"00000000",
		16#58a2# => X"00000000",
		16#58a3# => X"00000000",
		16#58a4# => X"00000000",
		16#58a5# => X"00000000",
		16#58a6# => X"00000000",
		16#58a7# => X"00000000",
		16#58a8# => X"00000000",
		16#58a9# => X"00000000",
		16#58aa# => X"00000000",
		16#58ab# => X"00000000",
		16#58ac# => X"00000000",
		16#58ad# => X"00000000",
		16#58ae# => X"00000000",
		16#58af# => X"00000000",
		16#58b0# => X"00000000",
		16#58b1# => X"00000000",
		16#58b2# => X"00000000",
		16#58b3# => X"00000000",
		16#58b4# => X"00000000",
		16#58b5# => X"00000000",
		16#58b6# => X"00000000",
		16#58b7# => X"00000000",
		16#58b8# => X"00000000",
		16#58b9# => X"00000000",
		16#58ba# => X"00000000",
		16#58bb# => X"00000000",
		16#58bc# => X"00000000",
		16#58bd# => X"00000000",
		16#58be# => X"00000000",
		16#58bf# => X"00000000",
		16#58c0# => X"00000000",
		16#58c1# => X"00000000",
		16#58c2# => X"00000000",
		16#58c3# => X"00000000",
		16#58c4# => X"00000000",
		16#58c5# => X"00000000",
		16#58c6# => X"00000000",
		16#58c7# => X"00000000",
		16#58c8# => X"00000000",
		16#58c9# => X"00000000",
		16#58ca# => X"00000000",
		16#58cb# => X"00000000",
		16#58cc# => X"00000000",
		16#58cd# => X"00000000",
		16#58ce# => X"00000000",
		16#58cf# => X"00000000",
		16#58d0# => X"00000000",
		16#58d1# => X"00000000",
		16#58d2# => X"00000000",
		16#58d3# => X"00000000",
		16#58d4# => X"00000000",
		16#58d5# => X"00000000",
		16#58d6# => X"00000000",
		16#58d7# => X"00000000",
		16#58d8# => X"00000000",
		16#58d9# => X"00000000",
		16#58da# => X"00000000",
		16#58db# => X"00000000",
		16#58dc# => X"00000000",
		16#58dd# => X"00000000",
		16#58de# => X"00000000",
		16#58df# => X"00000000",
		16#58e0# => X"00000000",
		16#58e1# => X"00000000",
		16#58e2# => X"00000000",
		16#58e3# => X"00000000",
		16#58e4# => X"00000000",
		16#58e5# => X"00000000",
		16#58e6# => X"00000000",
		16#58e7# => X"00000000",
		16#58e8# => X"00000000",
		16#58e9# => X"00000000",
		16#58ea# => X"00000000",
		16#58eb# => X"00000000",
		16#58ec# => X"00000000",
		16#58ed# => X"00000000",
		16#58ee# => X"00000000",
		16#58ef# => X"00000000",
		16#58f0# => X"00000000",
		16#58f1# => X"00000000",
		16#58f2# => X"00000000",
		16#58f3# => X"00000000",
		16#58f4# => X"00000000",
		16#58f5# => X"00000000",
		16#58f6# => X"00000000",
		16#58f7# => X"00000000",
		16#58f8# => X"00000000",
		16#58f9# => X"00000000",
		16#58fa# => X"00000000",
		16#58fb# => X"00000000",
		16#58fc# => X"00000000",
		16#58fd# => X"00000000",
		16#58fe# => X"00000000",
		16#58ff# => X"00000000",
		16#5900# => X"00000000",
		16#5901# => X"00000000",
		16#5902# => X"00000000",
		16#5903# => X"00000000",
		16#5904# => X"00000000",
		16#5905# => X"00000000",
		16#5906# => X"00000000",
		16#5907# => X"00000000",
		16#5908# => X"00000000",
		16#5909# => X"00000000",
		16#590a# => X"00000000",
		16#590b# => X"00000000",
		16#590c# => X"00000000",
		16#590d# => X"00000000",
		16#590e# => X"00000000",
		16#590f# => X"00000000",
		16#5910# => X"00000000",
		16#5911# => X"00000000",
		16#5912# => X"00000000",
		16#5913# => X"00000000",
		16#5914# => X"00000000",
		16#5915# => X"00000000",
		16#5916# => X"00000000",
		16#5917# => X"00000000",
		16#5918# => X"00000000",
		16#5919# => X"00000000",
		16#591a# => X"00000000",
		16#591b# => X"00000000",
		16#591c# => X"00000000",
		16#591d# => X"00000000",
		16#591e# => X"00000000",
		16#591f# => X"00000000",
		16#5920# => X"00000000",
		16#5921# => X"00000000",
		16#5922# => X"00000000",
		16#5923# => X"00000000",
		16#5924# => X"00000000",
		16#5925# => X"00000000",
		16#5926# => X"00000000",
		16#5927# => X"00000000",
		16#5928# => X"00000000",
		16#5929# => X"00000000",
		16#592a# => X"00000000",
		16#592b# => X"00000000",
		16#592c# => X"00000000",
		16#592d# => X"00000000",
		16#592e# => X"00000000",
		16#592f# => X"00000000",
		16#5930# => X"00000000",
		16#5931# => X"00000000",
		16#5932# => X"00000000",
		16#5933# => X"00000000",
		16#5934# => X"00000000",
		16#5935# => X"00000000",
		16#5936# => X"00000000",
		16#5937# => X"00000000",
		16#5938# => X"00000000",
		16#5939# => X"00000000",
		16#593a# => X"00000000",
		16#593b# => X"00000000",
		16#593c# => X"00000000",
		16#593d# => X"00000000",
		16#593e# => X"00000000",
		16#593f# => X"00000000",
		16#5940# => X"00000000",
		16#5941# => X"00000000",
		16#5942# => X"00000000",
		16#5943# => X"00000000",
		16#5944# => X"00000000",
		16#5945# => X"00000000",
		16#5946# => X"00000000",
		16#5947# => X"00000000",
		16#5948# => X"00000000",
		16#5949# => X"00000000",
		16#594a# => X"00000000",
		16#594b# => X"00000000",
		16#594c# => X"00000000",
		16#594d# => X"00000000",
		16#594e# => X"00000000",
		16#594f# => X"00000000",
		16#5950# => X"00000000",
		16#5951# => X"00000000",
		16#5952# => X"00000000",
		16#5953# => X"00000000",
		16#5954# => X"00000000",
		16#5955# => X"00000000",
		16#5956# => X"00000000",
		16#5957# => X"00000000",
		16#5958# => X"00000000",
		16#5959# => X"00000000",
		16#595a# => X"00000000",
		16#595b# => X"00000000",
		16#595c# => X"00000000",
		16#595d# => X"00000000",
		16#595e# => X"00000000",
		16#595f# => X"00000000",
		16#5960# => X"00000000",
		16#5961# => X"00000000",
		16#5962# => X"00000000",
		16#5963# => X"00000000",
		16#5964# => X"00000000",
		16#5965# => X"00000000",
		16#5966# => X"00000000",
		16#5967# => X"00000000",
		16#5968# => X"00000000",
		16#5969# => X"00000000",
		16#596a# => X"00000000",
		16#596b# => X"00000000",
		16#596c# => X"00000000",
		16#596d# => X"00000000",
		16#596e# => X"00000000",
		16#596f# => X"00000000",
		16#5970# => X"00000000",
		16#5971# => X"00000000",
		16#5972# => X"00000000",
		16#5973# => X"00000000",
		16#5974# => X"00000000",
		16#5975# => X"00000000",
		16#5976# => X"00000000",
		16#5977# => X"00000000",
		16#5978# => X"00000000",
		16#5979# => X"00000000",
		16#597a# => X"00000000",
		16#597b# => X"00000000",
		16#597c# => X"00000000",
		16#597d# => X"00000000",
		16#597e# => X"00000000",
		16#597f# => X"00000000",
		16#5980# => X"00000000",
		16#5981# => X"00000000",
		16#5982# => X"00000000",
		16#5983# => X"00000000",
		16#5984# => X"00000000",
		16#5985# => X"00000000",
		16#5986# => X"00000000",
		16#5987# => X"00000000",
		16#5988# => X"00000000",
		16#5989# => X"00000000",
		16#598a# => X"00000000",
		16#598b# => X"00000000",
		16#598c# => X"00000000",
		16#598d# => X"00000000",
		16#598e# => X"00000000",
		16#598f# => X"00000000",
		16#5990# => X"00000000",
		16#5991# => X"00000000",
		16#5992# => X"00000000",
		16#5993# => X"00000000",
		16#5994# => X"00000000",
		16#5995# => X"00000000",
		16#5996# => X"00000000",
		16#5997# => X"00000000",
		16#5998# => X"00000000",
		16#5999# => X"00000000",
		16#599a# => X"00000000",
		16#599b# => X"00000000",
		16#599c# => X"00000000",
		16#599d# => X"00000000",
		16#599e# => X"00000000",
		16#599f# => X"00000000",
		16#59a0# => X"00000000",
		16#59a1# => X"00000000",
		16#59a2# => X"00000000",
		16#59a3# => X"00000000",
		16#59a4# => X"00000000",
		16#59a5# => X"00000000",
		16#59a6# => X"00000000",
		16#59a7# => X"00000000",
		16#59a8# => X"00000000",
		16#59a9# => X"00000000",
		16#59aa# => X"00000000",
		16#59ab# => X"00000000",
		16#59ac# => X"00000000",
		16#59ad# => X"00000000",
		16#59ae# => X"00000000",
		16#59af# => X"00000000",
		16#59b0# => X"00000000",
		16#59b1# => X"00000000",
		16#59b2# => X"00000000",
		16#59b3# => X"00000000",
		16#59b4# => X"00000000",
		16#59b5# => X"00000000",
		16#59b6# => X"00000000",
		16#59b7# => X"00000000",
		16#59b8# => X"00000000",
		16#59b9# => X"00000000",
		16#59ba# => X"00000000",
		16#59bb# => X"00000000",
		16#59bc# => X"00000000",
		16#59bd# => X"00000000",
		16#59be# => X"00000000",
		16#59bf# => X"00000000",
		16#59c0# => X"00000000",
		16#59c1# => X"00000000",
		16#59c2# => X"00000000",
		16#59c3# => X"00000000",
		16#59c4# => X"00000000",
		16#59c5# => X"00000000",
		16#59c6# => X"00000000",
		16#59c7# => X"00000000",
		16#59c8# => X"00000000",
		16#59c9# => X"00000000",
		16#59ca# => X"00000000",
		16#59cb# => X"00000000",
		16#59cc# => X"00000000",
		16#59cd# => X"00000000",
		16#59ce# => X"00000000",
		16#59cf# => X"00000000",
		16#59d0# => X"00000000",
		16#59d1# => X"00000000",
		16#59d2# => X"00000000",
		16#59d3# => X"00000000",
		16#59d4# => X"00000000",
		16#59d5# => X"00000000",
		16#59d6# => X"00000000",
		16#59d7# => X"00000000",
		16#59d8# => X"00000000",
		16#59d9# => X"00000000",
		16#59da# => X"00000000",
		16#59db# => X"00000000",
		16#59dc# => X"00000000",
		16#59dd# => X"00000000",
		16#59de# => X"00000000",
		16#59df# => X"00000000",
		16#59e0# => X"00000000",
		16#59e1# => X"00000000",
		16#59e2# => X"00000000",
		16#59e3# => X"00000000",
		16#59e4# => X"00000000",
		16#59e5# => X"00000000",
		16#59e6# => X"00000000",
		16#59e7# => X"00000000",
		16#59e8# => X"00000000",
		16#59e9# => X"00000000",
		16#59ea# => X"00000000",
		16#59eb# => X"00000000",
		16#59ec# => X"00000000",
		16#59ed# => X"00000000",
		16#59ee# => X"00000000",
		16#59ef# => X"00000000",
		16#59f0# => X"00000000",
		16#59f1# => X"00000000",
		16#59f2# => X"00000000",
		16#59f3# => X"00000000",
		16#59f4# => X"00000000",
		16#59f5# => X"00000000",
		16#59f6# => X"00000000",
		16#59f7# => X"00000000",
		16#59f8# => X"00000000",
		16#59f9# => X"00000000",
		16#59fa# => X"00000000",
		16#59fb# => X"00000000",
		16#59fc# => X"00000000",
		16#59fd# => X"00000000",
		16#59fe# => X"00000000",
		16#59ff# => X"00000000",
		16#5a00# => X"00000000",
		16#5a01# => X"00000000",
		16#5a02# => X"00000000",
		16#5a03# => X"00000000",
		16#5a04# => X"00000000",
		16#5a05# => X"00000000",
		16#5a06# => X"00000000",
		16#5a07# => X"00000000",
		16#5a08# => X"00000000",
		16#5a09# => X"00000000",
		16#5a0a# => X"00000000",
		16#5a0b# => X"00000000",
		16#5a0c# => X"00000000",
		16#5a0d# => X"00000000",
		16#5a0e# => X"00000000",
		16#5a0f# => X"00000000",
		16#5a10# => X"00000000",
		16#5a11# => X"00000000",
		16#5a12# => X"00000000",
		16#5a13# => X"00000000",
		16#5a14# => X"00000000",
		16#5a15# => X"00000000",
		16#5a16# => X"00000000",
		16#5a17# => X"00000000",
		16#5a18# => X"00000000",
		16#5a19# => X"00000000",
		16#5a1a# => X"00000000",
		16#5a1b# => X"00000000",
		16#5a1c# => X"00000000",
		16#5a1d# => X"00000000",
		16#5a1e# => X"00000000",
		16#5a1f# => X"00000000",
		16#5a20# => X"00000000",
		16#5a21# => X"00000000",
		16#5a22# => X"00000000",
		16#5a23# => X"00000000",
		16#5a24# => X"00000000",
		16#5a25# => X"00000000",
		16#5a26# => X"00000000",
		16#5a27# => X"00000000",
		16#5a28# => X"00000000",
		16#5a29# => X"00000000",
		16#5a2a# => X"00000000",
		16#5a2b# => X"00000000",
		16#5a2c# => X"00000000",
		16#5a2d# => X"00000000",
		16#5a2e# => X"00000000",
		16#5a2f# => X"00000000",
		16#5a30# => X"00000000",
		16#5a31# => X"00000000",
		16#5a32# => X"00000000",
		16#5a33# => X"00000000",
		16#5a34# => X"00000000",
		16#5a35# => X"00000000",
		16#5a36# => X"00000000",
		16#5a37# => X"00000000",
		16#5a38# => X"00000000",
		16#5a39# => X"00000000",
		16#5a3a# => X"00000000",
		16#5a3b# => X"00000000",
		16#5a3c# => X"00000000",
		16#5a3d# => X"00000000",
		16#5a3e# => X"00000000",
		16#5a3f# => X"00000000",
		16#5a40# => X"00000000",
		16#5a41# => X"00000000",
		16#5a42# => X"00000000",
		16#5a43# => X"00000000",
		16#5a44# => X"00000000",
		16#5a45# => X"00000000",
		16#5a46# => X"00000000",
		16#5a47# => X"00000000",
		16#5a48# => X"00000000",
		16#5a49# => X"00000000",
		16#5a4a# => X"00000000",
		16#5a4b# => X"00000000",
		16#5a4c# => X"00000000",
		16#5a4d# => X"00000000",
		16#5a4e# => X"00000000",
		16#5a4f# => X"00000000",
		16#5a50# => X"00000000",
		16#5a51# => X"00000000",
		16#5a52# => X"00000000",
		16#5a53# => X"00000000",
		16#5a54# => X"00000000",
		16#5a55# => X"00000000",
		16#5a56# => X"00000000",
		16#5a57# => X"00000000",
		16#5a58# => X"00000000",
		16#5a59# => X"00000000",
		16#5a5a# => X"00000000",
		16#5a5b# => X"00000000",
		16#5a5c# => X"00000000",
		16#5a5d# => X"00000000",
		16#5a5e# => X"00000000",
		16#5a5f# => X"00000000",
		16#5a60# => X"00000000",
		16#5a61# => X"00000000",
		16#5a62# => X"00000000",
		16#5a63# => X"00000000",
		16#5a64# => X"00000000",
		16#5a65# => X"00000000",
		16#5a66# => X"00000000",
		16#5a67# => X"00000000",
		16#5a68# => X"00000000",
		16#5a69# => X"00000000",
		16#5a6a# => X"00000000",
		16#5a6b# => X"00000000",
		16#5a6c# => X"00000000",
		16#5a6d# => X"00000000",
		16#5a6e# => X"00000000",
		16#5a6f# => X"00000000",
		16#5a70# => X"00000000",
		16#5a71# => X"00000000",
		16#5a72# => X"00000000",
		16#5a73# => X"00000000",
		16#5a74# => X"00000000",
		16#5a75# => X"00000000",
		16#5a76# => X"00000000",
		16#5a77# => X"00000000",
		16#5a78# => X"00000000",
		16#5a79# => X"00000000",
		16#5a7a# => X"00000000",
		16#5a7b# => X"00000000",
		16#5a7c# => X"00000000",
		16#5a7d# => X"00000000",
		16#5a7e# => X"00000000",
		16#5a7f# => X"00000000",
		16#5a80# => X"00000000",
		16#5a81# => X"00000000",
		16#5a82# => X"00000000",
		16#5a83# => X"00000000",
		16#5a84# => X"00000000",
		16#5a85# => X"00000000",
		16#5a86# => X"00000000",
		16#5a87# => X"00000000",
		16#5a88# => X"00000000",
		16#5a89# => X"00000000",
		16#5a8a# => X"00000000",
		16#5a8b# => X"00000000",
		16#5a8c# => X"00000000",
		16#5a8d# => X"00000000",
		16#5a8e# => X"00000000",
		16#5a8f# => X"00000000",
		16#5a90# => X"00000000",
		16#5a91# => X"00000000",
		16#5a92# => X"00000000",
		16#5a93# => X"00000000",
		16#5a94# => X"00000000",
		16#5a95# => X"00000000",
		16#5a96# => X"00000000",
		16#5a97# => X"00000000",
		16#5a98# => X"00000000",
		16#5a99# => X"00000000",
		16#5a9a# => X"00000000",
		16#5a9b# => X"00000000",
		16#5a9c# => X"00000000",
		16#5a9d# => X"00000000",
		16#5a9e# => X"00000000",
		16#5a9f# => X"00000000",
		16#5aa0# => X"00000000",
		16#5aa1# => X"00000000",
		16#5aa2# => X"00000000",
		16#5aa3# => X"00000000",
		16#5aa4# => X"00000000",
		16#5aa5# => X"00000000",
		16#5aa6# => X"00000000",
		16#5aa7# => X"00000000",
		16#5aa8# => X"00000000",
		16#5aa9# => X"00000000",
		16#5aaa# => X"00000000",
		16#5aab# => X"00000000",
		16#5aac# => X"00000000",
		16#5aad# => X"00000000",
		16#5aae# => X"00000000",
		16#5aaf# => X"00000000",
		16#5ab0# => X"00000000",
		16#5ab1# => X"00000000",
		16#5ab2# => X"00000000",
		16#5ab3# => X"00000000",
		16#5ab4# => X"00000000",
		16#5ab5# => X"00000000",
		16#5ab6# => X"00000000",
		16#5ab7# => X"00000000",
		16#5ab8# => X"00000000",
		16#5ab9# => X"00000000",
		16#5aba# => X"00000000",
		16#5abb# => X"00000000",
		16#5abc# => X"00000000",
		16#5abd# => X"00000000",
		16#5abe# => X"00000000",
		16#5abf# => X"00000000",
		16#5ac0# => X"00000000",
		16#5ac1# => X"00000000",
		16#5ac2# => X"00000000",
		16#5ac3# => X"00000000",
		16#5ac4# => X"00000000",
		16#5ac5# => X"00000000",
		16#5ac6# => X"00000000",
		16#5ac7# => X"00000000",
		16#5ac8# => X"00000000",
		16#5ac9# => X"00000000",
		16#5aca# => X"00000000",
		16#5acb# => X"00000000",
		16#5acc# => X"00000000",
		16#5acd# => X"00000000",
		16#5ace# => X"00000000",
		16#5acf# => X"00000000",
		16#5ad0# => X"00000000",
		16#5ad1# => X"00000000",
		16#5ad2# => X"00000000",
		16#5ad3# => X"00000000",
		16#5ad4# => X"00000000",
		16#5ad5# => X"00000000",
		16#5ad6# => X"00000000",
		16#5ad7# => X"00000000",
		16#5ad8# => X"00000000",
		16#5ad9# => X"00000000",
		16#5ada# => X"00000000",
		16#5adb# => X"00000000",
		16#5adc# => X"00000000",
		16#5add# => X"00000000",
		16#5ade# => X"00000000",
		16#5adf# => X"00000000",
		16#5ae0# => X"00000000",
		16#5ae1# => X"00000000",
		16#5ae2# => X"00000000",
		16#5ae3# => X"00000000",
		16#5ae4# => X"00000000",
		16#5ae5# => X"00000000",
		16#5ae6# => X"00000000",
		16#5ae7# => X"00000000",
		16#5ae8# => X"00000000",
		16#5ae9# => X"00000000",
		16#5aea# => X"00000000",
		16#5aeb# => X"00000000",
		16#5aec# => X"00000000",
		16#5aed# => X"00000000",
		16#5aee# => X"00000000",
		16#5aef# => X"00000000",
		16#5af0# => X"00000000",
		16#5af1# => X"00000000",
		16#5af2# => X"00000000",
		16#5af3# => X"00000000",
		16#5af4# => X"00000000",
		16#5af5# => X"00000000",
		16#5af6# => X"00000000",
		16#5af7# => X"00000000",
		16#5af8# => X"00000000",
		16#5af9# => X"00000000",
		16#5afa# => X"00000000",
		16#5afb# => X"00000000",
		16#5afc# => X"00000000",
		16#5afd# => X"00000000",
		16#5afe# => X"00000000",
		16#5aff# => X"00000000",
		16#5b00# => X"00000000",
		16#5b01# => X"00000000",
		16#5b02# => X"00000000",
		16#5b03# => X"00000000",
		16#5b04# => X"00000000",
		16#5b05# => X"00000000",
		16#5b06# => X"00000000",
		16#5b07# => X"00000000",
		16#5b08# => X"00000000",
		16#5b09# => X"00000000",
		16#5b0a# => X"00000000",
		16#5b0b# => X"00000000",
		16#5b0c# => X"00000000",
		16#5b0d# => X"00000000",
		16#5b0e# => X"00000000",
		16#5b0f# => X"00000000",
		16#5b10# => X"00000000",
		16#5b11# => X"00000000",
		16#5b12# => X"00000000",
		16#5b13# => X"00000000",
		16#5b14# => X"00000000",
		16#5b15# => X"00000000",
		16#5b16# => X"00000000",
		16#5b17# => X"00000000",
		16#5b18# => X"00000000",
		16#5b19# => X"00000000",
		16#5b1a# => X"00000000",
		16#5b1b# => X"00000000",
		16#5b1c# => X"00000000",
		16#5b1d# => X"00000000",
		16#5b1e# => X"00000000",
		16#5b1f# => X"00000000",
		16#5b20# => X"00000000",
		16#5b21# => X"00000000",
		16#5b22# => X"00000000",
		16#5b23# => X"00000000",
		16#5b24# => X"00000000",
		16#5b25# => X"00000000",
		16#5b26# => X"00000000",
		16#5b27# => X"00000000",
		16#5b28# => X"00000000",
		16#5b29# => X"00000000",
		16#5b2a# => X"00000000",
		16#5b2b# => X"00000000",
		16#5b2c# => X"00000000",
		16#5b2d# => X"00000000",
		16#5b2e# => X"00000000",
		16#5b2f# => X"00000000",
		16#5b30# => X"00000000",
		16#5b31# => X"00000000",
		16#5b32# => X"00000000",
		16#5b33# => X"00000000",
		16#5b34# => X"00000000",
		16#5b35# => X"00000000",
		16#5b36# => X"00000000",
		16#5b37# => X"00000000",
		16#5b38# => X"00000000",
		16#5b39# => X"00000000",
		16#5b3a# => X"00000000",
		16#5b3b# => X"00000000",
		16#5b3c# => X"00000000",
		16#5b3d# => X"00000000",
		16#5b3e# => X"00000000",
		16#5b3f# => X"00000000",
		16#5b40# => X"00000000",
		16#5b41# => X"00000000",
		16#5b42# => X"00000000",
		16#5b43# => X"00000000",
		16#5b44# => X"00000000",
		16#5b45# => X"00000000",
		16#5b46# => X"00000000",
		16#5b47# => X"00000000",
		16#5b48# => X"00000000",
		16#5b49# => X"00000000",
		16#5b4a# => X"00000000",
		16#5b4b# => X"00000000",
		16#5b4c# => X"00000000",
		16#5b4d# => X"00000000",
		16#5b4e# => X"00000000",
		16#5b4f# => X"00000000",
		16#5b50# => X"00000000",
		16#5b51# => X"00000000",
		16#5b52# => X"00000000",
		16#5b53# => X"00000000",
		16#5b54# => X"00000000",
		16#5b55# => X"00000000",
		16#5b56# => X"00000000",
		16#5b57# => X"00000000",
		16#5b58# => X"00000000",
		16#5b59# => X"00000000",
		16#5b5a# => X"00000000",
		16#5b5b# => X"00000000",
		16#5b5c# => X"00000000",
		16#5b5d# => X"00000000",
		16#5b5e# => X"00000000",
		16#5b5f# => X"00000000",
		16#5b60# => X"00000000",
		16#5b61# => X"00000000",
		16#5b62# => X"00000000",
		16#5b63# => X"00000000",
		16#5b64# => X"00000000",
		16#5b65# => X"00000000",
		16#5b66# => X"00000000",
		16#5b67# => X"00000000",
		16#5b68# => X"00000000",
		16#5b69# => X"00000000",
		16#5b6a# => X"00000000",
		16#5b6b# => X"00000000",
		16#5b6c# => X"00000000",
		16#5b6d# => X"00000000",
		16#5b6e# => X"00000000",
		16#5b6f# => X"00000000",
		16#5b70# => X"00000000",
		16#5b71# => X"00000000",
		16#5b72# => X"00000000",
		16#5b73# => X"00000000",
		16#5b74# => X"00000000",
		16#5b75# => X"00000000",
		16#5b76# => X"00000000",
		16#5b77# => X"00000000",
		16#5b78# => X"00000000",
		16#5b79# => X"00000000",
		16#5b7a# => X"00000000",
		16#5b7b# => X"00000000",
		16#5b7c# => X"00000000",
		16#5b7d# => X"00000000",
		16#5b7e# => X"00000000",
		16#5b7f# => X"00000000",
		16#5b80# => X"00000000",
		16#5b81# => X"00000000",
		16#5b82# => X"00000000",
		16#5b83# => X"00000000",
		16#5b84# => X"00000000",
		16#5b85# => X"00000000",
		16#5b86# => X"00000000",
		16#5b87# => X"00000000",
		16#5b88# => X"00000000",
		16#5b89# => X"00000000",
		16#5b8a# => X"00000000",
		16#5b8b# => X"00000000",
		16#5b8c# => X"00000000",
		16#5b8d# => X"00000000",
		16#5b8e# => X"00000000",
		16#5b8f# => X"00000000",
		16#5b90# => X"00000000",
		16#5b91# => X"00000000",
		16#5b92# => X"00000000",
		16#5b93# => X"00000000",
		16#5b94# => X"00000000",
		16#5b95# => X"00000000",
		16#5b96# => X"00000000",
		16#5b97# => X"00000000",
		16#5b98# => X"00000000",
		16#5b99# => X"00000000",
		16#5b9a# => X"00000000",
		16#5b9b# => X"00000000",
		16#5b9c# => X"00000000",
		16#5b9d# => X"00000000",
		16#5b9e# => X"00000000",
		16#5b9f# => X"00000000",
		16#5ba0# => X"00000000",
		16#5ba1# => X"00000000",
		16#5ba2# => X"00000000",
		16#5ba3# => X"00000000",
		16#5ba4# => X"00000000",
		16#5ba5# => X"00000000",
		16#5ba6# => X"00000000",
		16#5ba7# => X"00000000",
		16#5ba8# => X"00000000",
		16#5ba9# => X"00000000",
		16#5baa# => X"00000000",
		16#5bab# => X"00000000",
		16#5bac# => X"00000000",
		16#5bad# => X"00000000",
		16#5bae# => X"00000000",
		16#5baf# => X"00000000",
		16#5bb0# => X"00000000",
		16#5bb1# => X"00000000",
		16#5bb2# => X"00000000",
		16#5bb3# => X"00000000",
		16#5bb4# => X"00000000",
		16#5bb5# => X"00000000",
		16#5bb6# => X"00000000",
		16#5bb7# => X"00000000",
		16#5bb8# => X"00000000",
		16#5bb9# => X"00000000",
		16#5bba# => X"00000000",
		16#5bbb# => X"00000000",
		16#5bbc# => X"00000000",
		16#5bbd# => X"00000000",
		16#5bbe# => X"00000000",
		16#5bbf# => X"00000000",
		16#5bc0# => X"00000000",
		16#5bc1# => X"00000000",
		16#5bc2# => X"00000000",
		16#5bc3# => X"00000000",
		16#5bc4# => X"00000000",
		16#5bc5# => X"00000000",
		16#5bc6# => X"00000000",
		16#5bc7# => X"00000000",
		16#5bc8# => X"00000000",
		16#5bc9# => X"00000000",
		16#5bca# => X"00000000",
		16#5bcb# => X"00000000",
		16#5bcc# => X"00000000",
		16#5bcd# => X"00000000",
		16#5bce# => X"00000000",
		16#5bcf# => X"00000000",
		16#5bd0# => X"00000000",
		16#5bd1# => X"00000000",
		16#5bd2# => X"00000000",
		16#5bd3# => X"00000000",
		16#5bd4# => X"00000000",
		16#5bd5# => X"00000000",
		16#5bd6# => X"00000000",
		16#5bd7# => X"00000000",
		16#5bd8# => X"00000000",
		16#5bd9# => X"00000000",
		16#5bda# => X"00000000",
		16#5bdb# => X"00000000",
		16#5bdc# => X"00000000",
		16#5bdd# => X"00000000",
		16#5bde# => X"00000000",
		16#5bdf# => X"00000000",
		16#5be0# => X"00000000",
		16#5be1# => X"00000000",
		16#5be2# => X"00000000",
		16#5be3# => X"00000000",
		16#5be4# => X"00000000",
		16#5be5# => X"00000000",
		16#5be6# => X"00000000",
		16#5be7# => X"00000000",
		16#5be8# => X"00000000",
		16#5be9# => X"00000000",
		16#5bea# => X"00000000",
		16#5beb# => X"00000000",
		16#5bec# => X"00000000",
		16#5bed# => X"00000000",
		16#5bee# => X"00000000",
		16#5bef# => X"00000000",
		16#5bf0# => X"00000000",
		16#5bf1# => X"00000000",
		16#5bf2# => X"00000000",
		16#5bf3# => X"00000000",
		16#5bf4# => X"00000000",
		16#5bf5# => X"00000000",
		16#5bf6# => X"00000000",
		16#5bf7# => X"00000000",
		16#5bf8# => X"00000000",
		16#5bf9# => X"00000000",
		16#5bfa# => X"00000000",
		16#5bfb# => X"00000000",
		16#5bfc# => X"00000000",
		16#5bfd# => X"00000000",
		16#5bfe# => X"00000000",
		16#5bff# => X"00000000",
		16#5c00# => X"00000000",
		16#5c01# => X"00000000",
		16#5c02# => X"00000000",
		16#5c03# => X"00000000",
		16#5c04# => X"00000000",
		16#5c05# => X"00000000",
		16#5c06# => X"00000000",
		16#5c07# => X"00000000",
		16#5c08# => X"00000000",
		16#5c09# => X"00000000",
		16#5c0a# => X"00000000",
		16#5c0b# => X"00000000",
		16#5c0c# => X"00000000",
		16#5c0d# => X"00000000",
		16#5c0e# => X"00000000",
		16#5c0f# => X"00000000",
		16#5c10# => X"00000000",
		16#5c11# => X"00000000",
		16#5c12# => X"00000000",
		16#5c13# => X"00000000",
		16#5c14# => X"00000000",
		16#5c15# => X"00000000",
		16#5c16# => X"00000000",
		16#5c17# => X"00000000",
		16#5c18# => X"00000000",
		16#5c19# => X"00000000",
		16#5c1a# => X"00000000",
		16#5c1b# => X"00000000",
		16#5c1c# => X"00000000",
		16#5c1d# => X"00000000",
		16#5c1e# => X"00000000",
		16#5c1f# => X"00000000",
		16#5c20# => X"00000000",
		16#5c21# => X"00000000",
		16#5c22# => X"00000000",
		16#5c23# => X"00000000",
		16#5c24# => X"00000000",
		16#5c25# => X"00000000",
		16#5c26# => X"00000000",
		16#5c27# => X"00000000",
		16#5c28# => X"00000000",
		16#5c29# => X"00000000",
		16#5c2a# => X"00000000",
		16#5c2b# => X"00000000",
		16#5c2c# => X"00000000",
		16#5c2d# => X"00000000",
		16#5c2e# => X"00000000",
		16#5c2f# => X"00000000",
		16#5c30# => X"00000000",
		16#5c31# => X"00000000",
		16#5c32# => X"00000000",
		16#5c33# => X"00000000",
		16#5c34# => X"00000000",
		16#5c35# => X"00000000",
		16#5c36# => X"00000000",
		16#5c37# => X"00000000",
		16#5c38# => X"00000000",
		16#5c39# => X"00000000",
		16#5c3a# => X"00000000",
		16#5c3b# => X"00000000",
		16#5c3c# => X"00000000",
		16#5c3d# => X"00000000",
		16#5c3e# => X"00000000",
		16#5c3f# => X"00000000",
		16#5c40# => X"00000000",
		16#5c41# => X"00000000",
		16#5c42# => X"00000000",
		16#5c43# => X"00000000",
		16#5c44# => X"00000000",
		16#5c45# => X"00000000",
		16#5c46# => X"00000000",
		16#5c47# => X"00000000",
		16#5c48# => X"00000000",
		16#5c49# => X"00000000",
		16#5c4a# => X"00000000",
		16#5c4b# => X"00000000",
		16#5c4c# => X"00000000",
		16#5c4d# => X"00000000",
		16#5c4e# => X"00000000",
		16#5c4f# => X"00000000",
		16#5c50# => X"00000000",
		16#5c51# => X"00000000",
		16#5c52# => X"00000000",
		16#5c53# => X"00000000",
		16#5c54# => X"00000000",
		16#5c55# => X"00000000",
		16#5c56# => X"00000000",
		16#5c57# => X"00000000",
		16#5c58# => X"00000000",
		16#5c59# => X"00000000",
		16#5c5a# => X"00000000",
		16#5c5b# => X"00000000",
		16#5c5c# => X"00000000",
		16#5c5d# => X"00000000",
		16#5c5e# => X"00000000",
		16#5c5f# => X"00000000",
		16#5c60# => X"00000000",
		16#5c61# => X"00000000",
		16#5c62# => X"00000000",
		16#5c63# => X"00000000",
		16#5c64# => X"00000000",
		16#5c65# => X"00000000",
		16#5c66# => X"00000000",
		16#5c67# => X"00000000",
		16#5c68# => X"00000000",
		16#5c69# => X"00000000",
		16#5c6a# => X"00000000",
		16#5c6b# => X"00000000",
		16#5c6c# => X"00000000",
		16#5c6d# => X"00000000",
		16#5c6e# => X"00000000",
		16#5c6f# => X"00000000",
		16#5c70# => X"00000000",
		16#5c71# => X"00000000",
		16#5c72# => X"00000000",
		16#5c73# => X"00000000",
		16#5c74# => X"00000000",
		16#5c75# => X"00000000",
		16#5c76# => X"00000000",
		16#5c77# => X"00000000",
		16#5c78# => X"00000000",
		16#5c79# => X"00000000",
		16#5c7a# => X"00000000",
		16#5c7b# => X"00000000",
		16#5c7c# => X"00000000",
		16#5c7d# => X"00000000",
		16#5c7e# => X"00000000",
		16#5c7f# => X"00000000",
		16#5c80# => X"00000000",
		16#5c81# => X"00000000",
		16#5c82# => X"00000000",
		16#5c83# => X"00000000",
		16#5c84# => X"00000000",
		16#5c85# => X"00000000",
		16#5c86# => X"00000000",
		16#5c87# => X"00000000",
		16#5c88# => X"00000000",
		16#5c89# => X"00000000",
		16#5c8a# => X"00000000",
		16#5c8b# => X"00000000",
		16#5c8c# => X"00000000",
		16#5c8d# => X"00000000",
		16#5c8e# => X"00000000",
		16#5c8f# => X"00000000",
		16#5c90# => X"00000000",
		16#5c91# => X"00000000",
		16#5c92# => X"00000000",
		16#5c93# => X"00000000",
		16#5c94# => X"00000000",
		16#5c95# => X"00000000",
		16#5c96# => X"00000000",
		16#5c97# => X"00000000",
		16#5c98# => X"00000000",
		16#5c99# => X"00000000",
		16#5c9a# => X"00000000",
		16#5c9b# => X"00000000",
		16#5c9c# => X"00000000",
		16#5c9d# => X"00000000",
		16#5c9e# => X"00000000",
		16#5c9f# => X"00000000",
		16#5ca0# => X"00000000",
		16#5ca1# => X"00000000",
		16#5ca2# => X"00000000",
		16#5ca3# => X"00000000",
		16#5ca4# => X"00000000",
		16#5ca5# => X"00000000",
		16#5ca6# => X"00000000",
		16#5ca7# => X"00000000",
		16#5ca8# => X"00000000",
		16#5ca9# => X"00000000",
		16#5caa# => X"00000000",
		16#5cab# => X"00000000",
		16#5cac# => X"00000000",
		16#5cad# => X"00000000",
		16#5cae# => X"00000000",
		16#5caf# => X"00000000",
		16#5cb0# => X"00000000",
		16#5cb1# => X"00000000",
		16#5cb2# => X"00000000",
		16#5cb3# => X"00000000",
		16#5cb4# => X"00000000",
		16#5cb5# => X"00000000",
		16#5cb6# => X"00000000",
		16#5cb7# => X"00000000",
		16#5cb8# => X"00000000",
		16#5cb9# => X"00000000",
		16#5cba# => X"00000000",
		16#5cbb# => X"00000000",
		16#5cbc# => X"00000000",
		16#5cbd# => X"00000000",
		16#5cbe# => X"00000000",
		16#5cbf# => X"00000000",
		16#5cc0# => X"00000000",
		16#5cc1# => X"00000000",
		16#5cc2# => X"00000000",
		16#5cc3# => X"00000000",
		16#5cc4# => X"00000000",
		16#5cc5# => X"00000000",
		16#5cc6# => X"00000000",
		16#5cc7# => X"00000000",
		16#5cc8# => X"00000000",
		16#5cc9# => X"00000000",
		16#5cca# => X"00000000",
		16#5ccb# => X"00000000",
		16#5ccc# => X"00000000",
		16#5ccd# => X"00000000",
		16#5cce# => X"00000000",
		16#5ccf# => X"00000000",
		16#5cd0# => X"00000000",
		16#5cd1# => X"00000000",
		16#5cd2# => X"00000000",
		16#5cd3# => X"00000000",
		16#5cd4# => X"00000000",
		16#5cd5# => X"00000000",
		16#5cd6# => X"00000000",
		16#5cd7# => X"00000000",
		16#5cd8# => X"00000000",
		16#5cd9# => X"00000000",
		16#5cda# => X"00000000",
		16#5cdb# => X"00000000",
		16#5cdc# => X"00000000",
		16#5cdd# => X"00000000",
		16#5cde# => X"00000000",
		16#5cdf# => X"00000000",
		16#5ce0# => X"00000000",
		16#5ce1# => X"00000000",
		16#5ce2# => X"00000000",
		16#5ce3# => X"00000000",
		16#5ce4# => X"00000000",
		16#5ce5# => X"00000000",
		16#5ce6# => X"00000000",
		16#5ce7# => X"00000000",
		16#5ce8# => X"00000000",
		16#5ce9# => X"00000000",
		16#5cea# => X"00000000",
		16#5ceb# => X"00000000",
		16#5cec# => X"00000000",
		16#5ced# => X"00000000",
		16#5cee# => X"00000000",
		16#5cef# => X"00000000",
		16#5cf0# => X"00000000",
		16#5cf1# => X"00000000",
		16#5cf2# => X"00000000",
		16#5cf3# => X"00000000",
		16#5cf4# => X"00000000",
		16#5cf5# => X"00000000",
		16#5cf6# => X"00000000",
		16#5cf7# => X"00000000",
		16#5cf8# => X"00000000",
		16#5cf9# => X"00000000",
		16#5cfa# => X"00000000",
		16#5cfb# => X"00000000",
		16#5cfc# => X"00000000",
		16#5cfd# => X"00000000",
		16#5cfe# => X"00000000",
		16#5cff# => X"00000000",
		16#5d00# => X"00000000",
		16#5d01# => X"00000000",
		16#5d02# => X"00000000",
		16#5d03# => X"00000000",
		16#5d04# => X"00000000",
		16#5d05# => X"00000000",
		16#5d06# => X"00000000",
		16#5d07# => X"00000000",
		16#5d08# => X"00000000",
		16#5d09# => X"00000000",
		16#5d0a# => X"00000000",
		16#5d0b# => X"00000000",
		16#5d0c# => X"00000000",
		16#5d0d# => X"00000000",
		16#5d0e# => X"00000000",
		16#5d0f# => X"00000000",
		16#5d10# => X"00000000",
		16#5d11# => X"00000000",
		16#5d12# => X"00000000",
		16#5d13# => X"00000000",
		16#5d14# => X"00000000",
		16#5d15# => X"00000000",
		16#5d16# => X"00000000",
		16#5d17# => X"00000000",
		16#5d18# => X"00000000",
		16#5d19# => X"00000000",
		16#5d1a# => X"00000000",
		16#5d1b# => X"00000000",
		16#5d1c# => X"00000000",
		16#5d1d# => X"00000000",
		16#5d1e# => X"00000000",
		16#5d1f# => X"00000000",
		16#5d20# => X"00000000",
		16#5d21# => X"00000000",
		16#5d22# => X"00000000",
		16#5d23# => X"00000000",
		16#5d24# => X"00000000",
		16#5d25# => X"00000000",
		16#5d26# => X"00000000",
		16#5d27# => X"00000000",
		16#5d28# => X"00000000",
		16#5d29# => X"00000000",
		16#5d2a# => X"00000000",
		16#5d2b# => X"00000000",
		16#5d2c# => X"00000000",
		16#5d2d# => X"00000000",
		16#5d2e# => X"00000000",
		16#5d2f# => X"00000000",
		16#5d30# => X"00000000",
		16#5d31# => X"00000000",
		16#5d32# => X"00000000",
		16#5d33# => X"00000000",
		16#5d34# => X"00000000",
		16#5d35# => X"00000000",
		16#5d36# => X"00000000",
		16#5d37# => X"00000000",
		16#5d38# => X"00000000",
		16#5d39# => X"00000000",
		16#5d3a# => X"00000000",
		16#5d3b# => X"00000000",
		16#5d3c# => X"00000000",
		16#5d3d# => X"00000000",
		16#5d3e# => X"00000000",
		16#5d3f# => X"00000000",
		16#5d40# => X"00000000",
		16#5d41# => X"00000000",
		16#5d42# => X"00000000",
		16#5d43# => X"00000000",
		16#5d44# => X"00000000",
		16#5d45# => X"00000000",
		16#5d46# => X"00000000",
		16#5d47# => X"00000000",
		16#5d48# => X"00000000",
		16#5d49# => X"00000000",
		16#5d4a# => X"00000000",
		16#5d4b# => X"00000000",
		16#5d4c# => X"00000000",
		16#5d4d# => X"00000000",
		16#5d4e# => X"00000000",
		16#5d4f# => X"00000000",
		16#5d50# => X"00000000",
		16#5d51# => X"00000000",
		16#5d52# => X"00000000",
		16#5d53# => X"00000000",
		16#5d54# => X"00000000",
		16#5d55# => X"00000000",
		16#5d56# => X"00000000",
		16#5d57# => X"00000000",
		16#5d58# => X"00000000",
		16#5d59# => X"00000000",
		16#5d5a# => X"00000000",
		16#5d5b# => X"00000000",
		16#5d5c# => X"00000000",
		16#5d5d# => X"00000000",
		16#5d5e# => X"00000000",
		16#5d5f# => X"00000000",
		16#5d60# => X"00000000",
		16#5d61# => X"00000000",
		16#5d62# => X"00000000",
		16#5d63# => X"00000000",
		16#5d64# => X"00000000",
		16#5d65# => X"00000000",
		16#5d66# => X"00000000",
		16#5d67# => X"00000000",
		16#5d68# => X"00000000",
		16#5d69# => X"00000000",
		16#5d6a# => X"00000000",
		16#5d6b# => X"00000000",
		16#5d6c# => X"00000000",
		16#5d6d# => X"00000000",
		16#5d6e# => X"00000000",
		16#5d6f# => X"00000000",
		16#5d70# => X"00000000",
		16#5d71# => X"00000000",
		16#5d72# => X"00000000",
		16#5d73# => X"00000000",
		16#5d74# => X"00000000",
		16#5d75# => X"00000000",
		16#5d76# => X"00000000",
		16#5d77# => X"00000000",
		16#5d78# => X"00000000",
		16#5d79# => X"00000000",
		16#5d7a# => X"00000000",
		16#5d7b# => X"00000000",
		16#5d7c# => X"00000000",
		16#5d7d# => X"00000000",
		16#5d7e# => X"00000000",
		16#5d7f# => X"00000000",
		16#5d80# => X"00000000",
		16#5d81# => X"00000000",
		16#5d82# => X"00000000",
		16#5d83# => X"00000000",
		16#5d84# => X"00000000",
		16#5d85# => X"00000000",
		16#5d86# => X"00000000",
		16#5d87# => X"00000000",
		16#5d88# => X"00000000",
		16#5d89# => X"00000000",
		16#5d8a# => X"00000000",
		16#5d8b# => X"00000000",
		16#5d8c# => X"00000000",
		16#5d8d# => X"00000000",
		16#5d8e# => X"00000000",
		16#5d8f# => X"00000000",
		16#5d90# => X"00000000",
		16#5d91# => X"00000000",
		16#5d92# => X"00000000",
		16#5d93# => X"00000000",
		16#5d94# => X"00000000",
		16#5d95# => X"00000000",
		16#5d96# => X"00000000",
		16#5d97# => X"00000000",
		16#5d98# => X"00000000",
		16#5d99# => X"00000000",
		16#5d9a# => X"00000000",
		16#5d9b# => X"00000000",
		16#5d9c# => X"00000000",
		16#5d9d# => X"00000000",
		16#5d9e# => X"00000000",
		16#5d9f# => X"00000000",
		16#5da0# => X"00000000",
		16#5da1# => X"00000000",
		16#5da2# => X"00000000",
		16#5da3# => X"00000000",
		16#5da4# => X"00000000",
		16#5da5# => X"00000000",
		16#5da6# => X"00000000",
		16#5da7# => X"00000000",
		16#5da8# => X"00000000",
		16#5da9# => X"00000000",
		16#5daa# => X"00000000",
		16#5dab# => X"00000000",
		16#5dac# => X"00000000",
		16#5dad# => X"00000000",
		16#5dae# => X"00000000",
		16#5daf# => X"00000000",
		16#5db0# => X"00000000",
		16#5db1# => X"00000000",
		16#5db2# => X"00000000",
		16#5db3# => X"00000000",
		16#5db4# => X"00000000",
		16#5db5# => X"00000000",
		16#5db6# => X"00000000",
		16#5db7# => X"00000000",
		16#5db8# => X"00000000",
		16#5db9# => X"00000000",
		16#5dba# => X"00000000",
		16#5dbb# => X"00000000",
		16#5dbc# => X"00000000",
		16#5dbd# => X"00000000",
		16#5dbe# => X"00000000",
		16#5dbf# => X"00000000",
		16#5dc0# => X"00000000",
		16#5dc1# => X"00000000",
		16#5dc2# => X"00000000",
		16#5dc3# => X"00000000",
		16#5dc4# => X"00000000",
		16#5dc5# => X"00000000",
		16#5dc6# => X"00000000",
		16#5dc7# => X"00000000",
		16#5dc8# => X"00000000",
		16#5dc9# => X"00000000",
		16#5dca# => X"00000000",
		16#5dcb# => X"00000000",
		16#5dcc# => X"00000000",
		16#5dcd# => X"00000000",
		16#5dce# => X"00000000",
		16#5dcf# => X"00000000",
		16#5dd0# => X"00000000",
		16#5dd1# => X"00000000",
		16#5dd2# => X"00000000",
		16#5dd3# => X"00000000",
		16#5dd4# => X"00000000",
		16#5dd5# => X"00000000",
		16#5dd6# => X"00000000",
		16#5dd7# => X"00000000",
		16#5dd8# => X"00000000",
		16#5dd9# => X"00000000",
		16#5dda# => X"00000000",
		16#5ddb# => X"00000000",
		16#5ddc# => X"00000000",
		16#5ddd# => X"00000000",
		16#5dde# => X"00000000",
		16#5ddf# => X"00000000",
		16#5de0# => X"00000000",
		16#5de1# => X"00000000",
		16#5de2# => X"00000000",
		16#5de3# => X"00000000",
		16#5de4# => X"00000000",
		16#5de5# => X"00000000",
		16#5de6# => X"00000000",
		16#5de7# => X"00000000",
		16#5de8# => X"00000000",
		16#5de9# => X"00000000",
		16#5dea# => X"00000000",
		16#5deb# => X"00000000",
		16#5dec# => X"00000000",
		16#5ded# => X"00000000",
		16#5dee# => X"00000000",
		16#5def# => X"00000000",
		16#5df0# => X"00000000",
		16#5df1# => X"00000000",
		16#5df2# => X"00000000",
		16#5df3# => X"00000000",
		16#5df4# => X"00000000",
		16#5df5# => X"00000000",
		16#5df6# => X"00000000",
		16#5df7# => X"00000000",
		16#5df8# => X"00000000",
		16#5df9# => X"00000000",
		16#5dfa# => X"00000000",
		16#5dfb# => X"00000000",
		16#5dfc# => X"00000000",
		16#5dfd# => X"00000000",
		16#5dfe# => X"00000000",
		16#5dff# => X"00000000",
		16#5e00# => X"00000000",
		16#5e01# => X"00000000",
		16#5e02# => X"00000000",
		16#5e03# => X"00000000",
		16#5e04# => X"00000000",
		16#5e05# => X"00000000",
		16#5e06# => X"00000000",
		16#5e07# => X"00000000",
		16#5e08# => X"00000000",
		16#5e09# => X"00000000",
		16#5e0a# => X"00000000",
		16#5e0b# => X"00000000",
		16#5e0c# => X"00000000",
		16#5e0d# => X"00000000",
		16#5e0e# => X"00000000",
		16#5e0f# => X"00000000",
		16#5e10# => X"00000000",
		16#5e11# => X"00000000",
		16#5e12# => X"00000000",
		16#5e13# => X"00000000",
		16#5e14# => X"00000000",
		16#5e15# => X"00000000",
		16#5e16# => X"00000000",
		16#5e17# => X"00000000",
		16#5e18# => X"00000000",
		16#5e19# => X"00000000",
		16#5e1a# => X"00000000",
		16#5e1b# => X"00000000",
		16#5e1c# => X"00000000",
		16#5e1d# => X"00000000",
		16#5e1e# => X"00000000",
		16#5e1f# => X"00000000",
		16#5e20# => X"00000000",
		16#5e21# => X"00000000",
		16#5e22# => X"00000000",
		16#5e23# => X"00000000",
		16#5e24# => X"00000000",
		16#5e25# => X"00000000",
		16#5e26# => X"00000000",
		16#5e27# => X"00000000",
		16#5e28# => X"00000000",
		16#5e29# => X"00000000",
		16#5e2a# => X"00000000",
		16#5e2b# => X"00000000",
		16#5e2c# => X"00000000",
		16#5e2d# => X"00000000",
		16#5e2e# => X"00000000",
		16#5e2f# => X"00000000",
		16#5e30# => X"00000000",
		16#5e31# => X"00000000",
		16#5e32# => X"00000000",
		16#5e33# => X"00000000",
		16#5e34# => X"00000000",
		16#5e35# => X"00000000",
		16#5e36# => X"00000000",
		16#5e37# => X"00000000",
		16#5e38# => X"00000000",
		16#5e39# => X"00000000",
		16#5e3a# => X"00000000",
		16#5e3b# => X"00000000",
		16#5e3c# => X"00000000",
		16#5e3d# => X"00000000",
		16#5e3e# => X"00000000",
		16#5e3f# => X"00000000",
		16#5e40# => X"00000000",
		16#5e41# => X"00000000",
		16#5e42# => X"00000000",
		16#5e43# => X"00000000",
		16#5e44# => X"00000000",
		16#5e45# => X"00000000",
		16#5e46# => X"00000000",
		16#5e47# => X"00000000",
		16#5e48# => X"00000000",
		16#5e49# => X"00000000",
		16#5e4a# => X"00000000",
		16#5e4b# => X"00000000",
		16#5e4c# => X"00000000",
		16#5e4d# => X"00000000",
		16#5e4e# => X"00000000",
		16#5e4f# => X"00000000",
		16#5e50# => X"00000000",
		16#5e51# => X"00000000",
		16#5e52# => X"00000000",
		16#5e53# => X"00000000",
		16#5e54# => X"00000000",
		16#5e55# => X"00000000",
		16#5e56# => X"00000000",
		16#5e57# => X"00000000",
		16#5e58# => X"00000000",
		16#5e59# => X"00000000",
		16#5e5a# => X"00000000",
		16#5e5b# => X"00000000",
		16#5e5c# => X"00000000",
		16#5e5d# => X"00000000",
		16#5e5e# => X"00000000",
		16#5e5f# => X"00000000",
		16#5e60# => X"00000000",
		16#5e61# => X"00000000",
		16#5e62# => X"00000000",
		16#5e63# => X"00000000",
		16#5e64# => X"00000000",
		16#5e65# => X"00000000",
		16#5e66# => X"00000000",
		16#5e67# => X"00000000",
		16#5e68# => X"00000000",
		16#5e69# => X"00000000",
		16#5e6a# => X"00000000",
		16#5e6b# => X"00000000",
		16#5e6c# => X"00000000",
		16#5e6d# => X"00000000",
		16#5e6e# => X"00000000",
		16#5e6f# => X"00000000",
		16#5e70# => X"00000000",
		16#5e71# => X"00000000",
		16#5e72# => X"00000000",
		16#5e73# => X"00000000",
		16#5e74# => X"00000000",
		16#5e75# => X"00000000",
		16#5e76# => X"00000000",
		16#5e77# => X"00000000",
		16#5e78# => X"00000000",
		16#5e79# => X"00000000",
		16#5e7a# => X"00000000",
		16#5e7b# => X"00000000",
		16#5e7c# => X"00000000",
		16#5e7d# => X"00000000",
		16#5e7e# => X"00000000",
		16#5e7f# => X"00000000",
		16#5e80# => X"00000000",
		16#5e81# => X"00000000",
		16#5e82# => X"00000000",
		16#5e83# => X"00000000",
		16#5e84# => X"00000000",
		16#5e85# => X"00000000",
		16#5e86# => X"00000000",
		16#5e87# => X"00000000",
		16#5e88# => X"00000000",
		16#5e89# => X"00000000",
		16#5e8a# => X"00000000",
		16#5e8b# => X"00000000",
		16#5e8c# => X"00000000",
		16#5e8d# => X"00000000",
		16#5e8e# => X"00000000",
		16#5e8f# => X"00000000",
		16#5e90# => X"00000000",
		16#5e91# => X"00000000",
		16#5e92# => X"00000000",
		16#5e93# => X"00000000",
		16#5e94# => X"00000000",
		16#5e95# => X"00000000",
		16#5e96# => X"00000000",
		16#5e97# => X"00000000",
		16#5e98# => X"00000000",
		16#5e99# => X"00000000",
		16#5e9a# => X"00000000",
		16#5e9b# => X"00000000",
		16#5e9c# => X"00000000",
		16#5e9d# => X"00000000",
		16#5e9e# => X"00000000",
		16#5e9f# => X"00000000",
		16#5ea0# => X"00000000",
		16#5ea1# => X"00000000",
		16#5ea2# => X"00000000",
		16#5ea3# => X"00000000",
		16#5ea4# => X"00000000",
		16#5ea5# => X"00000000",
		16#5ea6# => X"00000000",
		16#5ea7# => X"00000000",
		16#5ea8# => X"00000000",
		16#5ea9# => X"00000000",
		16#5eaa# => X"00000000",
		16#5eab# => X"00000000",
		16#5eac# => X"00000000",
		16#5ead# => X"00000000",
		16#5eae# => X"00000000",
		others => X"00000000"
	);

end package;