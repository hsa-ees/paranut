library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.types.all;

package prog_mem is

	constant PROG_SIZE : integer := 10068;

	constant PROG_DATA : mem_type(0 to PROG_SIZE/4-1) := (
		16#0000# => X"00000000",
		16#0001# => X"00000000",
		16#0002# => X"00000000",
		16#0003# => X"00000000",
		16#0004# => X"00000000",
		16#0005# => X"00000000",
		16#0006# => X"00000000",
		16#0007# => X"00000000",
		16#0008# => X"00000000",
		16#0009# => X"00000000",
		16#000a# => X"00000000",
		16#000b# => X"00000000",
		16#000c# => X"00000000",
		16#000d# => X"00000000",
		16#000e# => X"00000000",
		16#000f# => X"00000000",
		16#0010# => X"00000000",
		16#0011# => X"00000000",
		16#0012# => X"00000000",
		16#0013# => X"00000000",
		16#0014# => X"00000000",
		16#0015# => X"00000000",
		16#0016# => X"00000000",
		16#0017# => X"00000000",
		16#0018# => X"00000000",
		16#0019# => X"00000000",
		16#001a# => X"00000000",
		16#001b# => X"00000000",
		16#001c# => X"00000000",
		16#001d# => X"00000000",
		16#001e# => X"00000000",
		16#001f# => X"00000000",
		16#0020# => X"00000000",
		16#0021# => X"00000000",
		16#0022# => X"00000000",
		16#0023# => X"00000000",
		16#0024# => X"00000000",
		16#0025# => X"00000000",
		16#0026# => X"00000000",
		16#0027# => X"00000000",
		16#0028# => X"00000000",
		16#0029# => X"00000000",
		16#002a# => X"00000000",
		16#002b# => X"00000000",
		16#002c# => X"00000000",
		16#002d# => X"00000000",
		16#002e# => X"00000000",
		16#002f# => X"00000000",
		16#0030# => X"00000000",
		16#0031# => X"00000000",
		16#0032# => X"00000000",
		16#0033# => X"00000000",
		16#0034# => X"00000000",
		16#0035# => X"00000000",
		16#0036# => X"00000000",
		16#0037# => X"00000000",
		16#0038# => X"00000000",
		16#0039# => X"00000000",
		16#003a# => X"00000000",
		16#003b# => X"00000000",
		16#003c# => X"00000000",
		16#003d# => X"00000000",
		16#003e# => X"00000000",
		16#003f# => X"00000000",
		16#0040# => X"000007c0",
		16#0041# => X"15000000",
		16#0042# => X"00000000",
		16#0043# => X"00000000",
		16#0044# => X"00000000",
		16#0045# => X"00000000",
		16#0046# => X"00000000",
		16#0047# => X"00000000",
		16#0048# => X"00000000",
		16#0049# => X"00000000",
		16#004a# => X"00000000",
		16#004b# => X"00000000",
		16#004c# => X"00000000",
		16#004d# => X"00000000",
		16#004e# => X"00000000",
		16#004f# => X"00000000",
		16#0050# => X"00000000",
		16#0051# => X"00000000",
		16#0052# => X"00000000",
		16#0053# => X"00000000",
		16#0054# => X"00000000",
		16#0055# => X"00000000",
		16#0056# => X"00000000",
		16#0057# => X"00000000",
		16#0058# => X"00000000",
		16#0059# => X"00000000",
		16#005a# => X"00000000",
		16#005b# => X"00000000",
		16#005c# => X"00000000",
		16#005d# => X"00000000",
		16#005e# => X"00000000",
		16#005f# => X"00000000",
		16#0060# => X"00000000",
		16#0061# => X"00000000",
		16#0062# => X"00000000",
		16#0063# => X"00000000",
		16#0064# => X"00000000",
		16#0065# => X"00000000",
		16#0066# => X"00000000",
		16#0067# => X"00000000",
		16#0068# => X"00000000",
		16#0069# => X"00000000",
		16#006a# => X"00000000",
		16#006b# => X"00000000",
		16#006c# => X"00000000",
		16#006d# => X"00000000",
		16#006e# => X"00000000",
		16#006f# => X"00000000",
		16#0070# => X"00000000",
		16#0071# => X"00000000",
		16#0072# => X"00000000",
		16#0073# => X"00000000",
		16#0074# => X"00000000",
		16#0075# => X"00000000",
		16#0076# => X"00000000",
		16#0077# => X"00000000",
		16#0078# => X"00000000",
		16#0079# => X"00000000",
		16#007a# => X"00000000",
		16#007b# => X"00000000",
		16#007c# => X"00000000",
		16#007d# => X"00000000",
		16#007e# => X"00000000",
		16#007f# => X"00000000",
		16#0080# => X"00000000",
		16#0081# => X"00000000",
		16#0082# => X"00000000",
		16#0083# => X"00000000",
		16#0084# => X"00000000",
		16#0085# => X"00000000",
		16#0086# => X"00000000",
		16#0087# => X"00000000",
		16#0088# => X"00000000",
		16#0089# => X"00000000",
		16#008a# => X"00000000",
		16#008b# => X"00000000",
		16#008c# => X"00000000",
		16#008d# => X"00000000",
		16#008e# => X"00000000",
		16#008f# => X"00000000",
		16#0090# => X"00000000",
		16#0091# => X"00000000",
		16#0092# => X"00000000",
		16#0093# => X"00000000",
		16#0094# => X"00000000",
		16#0095# => X"00000000",
		16#0096# => X"00000000",
		16#0097# => X"00000000",
		16#0098# => X"00000000",
		16#0099# => X"00000000",
		16#009a# => X"00000000",
		16#009b# => X"00000000",
		16#009c# => X"00000000",
		16#009d# => X"00000000",
		16#009e# => X"00000000",
		16#009f# => X"00000000",
		16#00a0# => X"00000000",
		16#00a1# => X"00000000",
		16#00a2# => X"00000000",
		16#00a3# => X"00000000",
		16#00a4# => X"00000000",
		16#00a5# => X"00000000",
		16#00a6# => X"00000000",
		16#00a7# => X"00000000",
		16#00a8# => X"00000000",
		16#00a9# => X"00000000",
		16#00aa# => X"00000000",
		16#00ab# => X"00000000",
		16#00ac# => X"00000000",
		16#00ad# => X"00000000",
		16#00ae# => X"00000000",
		16#00af# => X"00000000",
		16#00b0# => X"00000000",
		16#00b1# => X"00000000",
		16#00b2# => X"00000000",
		16#00b3# => X"00000000",
		16#00b4# => X"00000000",
		16#00b5# => X"00000000",
		16#00b6# => X"00000000",
		16#00b7# => X"00000000",
		16#00b8# => X"00000000",
		16#00b9# => X"00000000",
		16#00ba# => X"00000000",
		16#00bb# => X"00000000",
		16#00bc# => X"00000000",
		16#00bd# => X"00000000",
		16#00be# => X"00000000",
		16#00bf# => X"00000000",
		16#00c0# => X"00000000",
		16#00c1# => X"00000000",
		16#00c2# => X"00000000",
		16#00c3# => X"00000000",
		16#00c4# => X"00000000",
		16#00c5# => X"00000000",
		16#00c6# => X"00000000",
		16#00c7# => X"00000000",
		16#00c8# => X"00000000",
		16#00c9# => X"00000000",
		16#00ca# => X"00000000",
		16#00cb# => X"00000000",
		16#00cc# => X"00000000",
		16#00cd# => X"00000000",
		16#00ce# => X"00000000",
		16#00cf# => X"00000000",
		16#00d0# => X"00000000",
		16#00d1# => X"00000000",
		16#00d2# => X"00000000",
		16#00d3# => X"00000000",
		16#00d4# => X"00000000",
		16#00d5# => X"00000000",
		16#00d6# => X"00000000",
		16#00d7# => X"00000000",
		16#00d8# => X"00000000",
		16#00d9# => X"00000000",
		16#00da# => X"00000000",
		16#00db# => X"00000000",
		16#00dc# => X"00000000",
		16#00dd# => X"00000000",
		16#00de# => X"00000000",
		16#00df# => X"00000000",
		16#00e0# => X"00000000",
		16#00e1# => X"00000000",
		16#00e2# => X"00000000",
		16#00e3# => X"00000000",
		16#00e4# => X"00000000",
		16#00e5# => X"00000000",
		16#00e6# => X"00000000",
		16#00e7# => X"00000000",
		16#00e8# => X"00000000",
		16#00e9# => X"00000000",
		16#00ea# => X"00000000",
		16#00eb# => X"00000000",
		16#00ec# => X"00000000",
		16#00ed# => X"00000000",
		16#00ee# => X"00000000",
		16#00ef# => X"00000000",
		16#00f0# => X"00000000",
		16#00f1# => X"00000000",
		16#00f2# => X"00000000",
		16#00f3# => X"00000000",
		16#00f4# => X"00000000",
		16#00f5# => X"00000000",
		16#00f6# => X"00000000",
		16#00f7# => X"00000000",
		16#00f8# => X"00000000",
		16#00f9# => X"00000000",
		16#00fa# => X"00000000",
		16#00fb# => X"00000000",
		16#00fc# => X"00000000",
		16#00fd# => X"00000000",
		16#00fe# => X"00000000",
		16#00ff# => X"00000000",
		16#0100# => X"00000000",
		16#0101# => X"00000000",
		16#0102# => X"00000000",
		16#0103# => X"00000000",
		16#0104# => X"00000000",
		16#0105# => X"00000000",
		16#0106# => X"00000000",
		16#0107# => X"00000000",
		16#0108# => X"00000000",
		16#0109# => X"00000000",
		16#010a# => X"00000000",
		16#010b# => X"00000000",
		16#010c# => X"00000000",
		16#010d# => X"00000000",
		16#010e# => X"00000000",
		16#010f# => X"00000000",
		16#0110# => X"00000000",
		16#0111# => X"00000000",
		16#0112# => X"00000000",
		16#0113# => X"00000000",
		16#0114# => X"00000000",
		16#0115# => X"00000000",
		16#0116# => X"00000000",
		16#0117# => X"00000000",
		16#0118# => X"00000000",
		16#0119# => X"00000000",
		16#011a# => X"00000000",
		16#011b# => X"00000000",
		16#011c# => X"00000000",
		16#011d# => X"00000000",
		16#011e# => X"00000000",
		16#011f# => X"00000000",
		16#0120# => X"00000000",
		16#0121# => X"00000000",
		16#0122# => X"00000000",
		16#0123# => X"00000000",
		16#0124# => X"00000000",
		16#0125# => X"00000000",
		16#0126# => X"00000000",
		16#0127# => X"00000000",
		16#0128# => X"00000000",
		16#0129# => X"00000000",
		16#012a# => X"00000000",
		16#012b# => X"00000000",
		16#012c# => X"00000000",
		16#012d# => X"00000000",
		16#012e# => X"00000000",
		16#012f# => X"00000000",
		16#0130# => X"00000000",
		16#0131# => X"00000000",
		16#0132# => X"00000000",
		16#0133# => X"00000000",
		16#0134# => X"00000000",
		16#0135# => X"00000000",
		16#0136# => X"00000000",
		16#0137# => X"00000000",
		16#0138# => X"00000000",
		16#0139# => X"00000000",
		16#013a# => X"00000000",
		16#013b# => X"00000000",
		16#013c# => X"00000000",
		16#013d# => X"00000000",
		16#013e# => X"00000000",
		16#013f# => X"00000000",
		16#0140# => X"00000000",
		16#0141# => X"00000000",
		16#0142# => X"00000000",
		16#0143# => X"00000000",
		16#0144# => X"00000000",
		16#0145# => X"00000000",
		16#0146# => X"00000000",
		16#0147# => X"00000000",
		16#0148# => X"00000000",
		16#0149# => X"00000000",
		16#014a# => X"00000000",
		16#014b# => X"00000000",
		16#014c# => X"00000000",
		16#014d# => X"00000000",
		16#014e# => X"00000000",
		16#014f# => X"00000000",
		16#0150# => X"00000000",
		16#0151# => X"00000000",
		16#0152# => X"00000000",
		16#0153# => X"00000000",
		16#0154# => X"00000000",
		16#0155# => X"00000000",
		16#0156# => X"00000000",
		16#0157# => X"00000000",
		16#0158# => X"00000000",
		16#0159# => X"00000000",
		16#015a# => X"00000000",
		16#015b# => X"00000000",
		16#015c# => X"00000000",
		16#015d# => X"00000000",
		16#015e# => X"00000000",
		16#015f# => X"00000000",
		16#0160# => X"00000000",
		16#0161# => X"00000000",
		16#0162# => X"00000000",
		16#0163# => X"00000000",
		16#0164# => X"00000000",
		16#0165# => X"00000000",
		16#0166# => X"00000000",
		16#0167# => X"00000000",
		16#0168# => X"00000000",
		16#0169# => X"00000000",
		16#016a# => X"00000000",
		16#016b# => X"00000000",
		16#016c# => X"00000000",
		16#016d# => X"00000000",
		16#016e# => X"00000000",
		16#016f# => X"00000000",
		16#0170# => X"00000000",
		16#0171# => X"00000000",
		16#0172# => X"00000000",
		16#0173# => X"00000000",
		16#0174# => X"00000000",
		16#0175# => X"00000000",
		16#0176# => X"00000000",
		16#0177# => X"00000000",
		16#0178# => X"00000000",
		16#0179# => X"00000000",
		16#017a# => X"00000000",
		16#017b# => X"00000000",
		16#017c# => X"00000000",
		16#017d# => X"00000000",
		16#017e# => X"00000000",
		16#017f# => X"00000000",
		16#0180# => X"18201500",
		16#0181# => X"d4800824",
		16#0182# => X"24000000",
		16#0183# => X"00000000",
		16#0184# => X"00000000",
		16#0185# => X"00000000",
		16#0186# => X"00000000",
		16#0187# => X"00000000",
		16#0188# => X"00000000",
		16#0189# => X"00000000",
		16#018a# => X"00000000",
		16#018b# => X"00000000",
		16#018c# => X"00000000",
		16#018d# => X"00000000",
		16#018e# => X"00000000",
		16#018f# => X"00000000",
		16#0190# => X"00000000",
		16#0191# => X"00000000",
		16#0192# => X"00000000",
		16#0193# => X"00000000",
		16#0194# => X"00000000",
		16#0195# => X"00000000",
		16#0196# => X"00000000",
		16#0197# => X"00000000",
		16#0198# => X"00000000",
		16#0199# => X"00000000",
		16#019a# => X"00000000",
		16#019b# => X"00000000",
		16#019c# => X"00000000",
		16#019d# => X"00000000",
		16#019e# => X"00000000",
		16#019f# => X"00000000",
		16#01a0# => X"00000000",
		16#01a1# => X"00000000",
		16#01a2# => X"00000000",
		16#01a3# => X"00000000",
		16#01a4# => X"00000000",
		16#01a5# => X"00000000",
		16#01a6# => X"00000000",
		16#01a7# => X"00000000",
		16#01a8# => X"00000000",
		16#01a9# => X"00000000",
		16#01aa# => X"00000000",
		16#01ab# => X"00000000",
		16#01ac# => X"00000000",
		16#01ad# => X"00000000",
		16#01ae# => X"00000000",
		16#01af# => X"00000000",
		16#01b0# => X"00000000",
		16#01b1# => X"00000000",
		16#01b2# => X"00000000",
		16#01b3# => X"00000000",
		16#01b4# => X"00000000",
		16#01b5# => X"00000000",
		16#01b6# => X"00000000",
		16#01b7# => X"00000000",
		16#01b8# => X"00000000",
		16#01b9# => X"00000000",
		16#01ba# => X"00000000",
		16#01bb# => X"00000000",
		16#01bc# => X"00000000",
		16#01bd# => X"00000000",
		16#01be# => X"00000000",
		16#01bf# => X"00000000",
		16#01c0# => X"18201500",
		16#01c1# => X"d480082c",
		16#01c2# => X"24000000",
		16#01c3# => X"00000000",
		16#01c4# => X"00000000",
		16#01c5# => X"00000000",
		16#01c6# => X"00000000",
		16#01c7# => X"00000000",
		16#01c8# => X"00000000",
		16#01c9# => X"00000000",
		16#01ca# => X"00000000",
		16#01cb# => X"00000000",
		16#01cc# => X"00000000",
		16#01cd# => X"00000000",
		16#01ce# => X"00000000",
		16#01cf# => X"00000000",
		16#01d0# => X"00000000",
		16#01d1# => X"00000000",
		16#01d2# => X"00000000",
		16#01d3# => X"00000000",
		16#01d4# => X"00000000",
		16#01d5# => X"00000000",
		16#01d6# => X"00000000",
		16#01d7# => X"00000000",
		16#01d8# => X"00000000",
		16#01d9# => X"00000000",
		16#01da# => X"00000000",
		16#01db# => X"00000000",
		16#01dc# => X"00000000",
		16#01dd# => X"00000000",
		16#01de# => X"00000000",
		16#01df# => X"00000000",
		16#01e0# => X"00000000",
		16#01e1# => X"00000000",
		16#01e2# => X"00000000",
		16#01e3# => X"00000000",
		16#01e4# => X"00000000",
		16#01e5# => X"00000000",
		16#01e6# => X"00000000",
		16#01e7# => X"00000000",
		16#01e8# => X"00000000",
		16#01e9# => X"00000000",
		16#01ea# => X"00000000",
		16#01eb# => X"00000000",
		16#01ec# => X"00000000",
		16#01ed# => X"00000000",
		16#01ee# => X"00000000",
		16#01ef# => X"00000000",
		16#01f0# => X"00000000",
		16#01f1# => X"00000000",
		16#01f2# => X"00000000",
		16#01f3# => X"00000000",
		16#01f4# => X"00000000",
		16#01f5# => X"00000000",
		16#01f6# => X"00000000",
		16#01f7# => X"00000000",
		16#01f8# => X"00000000",
		16#01f9# => X"00000000",
		16#01fa# => X"00000000",
		16#01fb# => X"00000000",
		16#01fc# => X"00000000",
		16#01fd# => X"00000000",
		16#01fe# => X"00000000",
		16#01ff# => X"00000000",
		16#0200# => X"00000000",
		16#0201# => X"00000000",
		16#0202# => X"00000000",
		16#0203# => X"00000000",
		16#0204# => X"00000000",
		16#0205# => X"00000000",
		16#0206# => X"00000000",
		16#0207# => X"00000000",
		16#0208# => X"00000000",
		16#0209# => X"00000000",
		16#020a# => X"00000000",
		16#020b# => X"00000000",
		16#020c# => X"00000000",
		16#020d# => X"00000000",
		16#020e# => X"00000000",
		16#020f# => X"00000000",
		16#0210# => X"00000000",
		16#0211# => X"00000000",
		16#0212# => X"00000000",
		16#0213# => X"00000000",
		16#0214# => X"00000000",
		16#0215# => X"00000000",
		16#0216# => X"00000000",
		16#0217# => X"00000000",
		16#0218# => X"00000000",
		16#0219# => X"00000000",
		16#021a# => X"00000000",
		16#021b# => X"00000000",
		16#021c# => X"00000000",
		16#021d# => X"00000000",
		16#021e# => X"00000000",
		16#021f# => X"00000000",
		16#0220# => X"00000000",
		16#0221# => X"00000000",
		16#0222# => X"00000000",
		16#0223# => X"00000000",
		16#0224# => X"00000000",
		16#0225# => X"00000000",
		16#0226# => X"00000000",
		16#0227# => X"00000000",
		16#0228# => X"00000000",
		16#0229# => X"00000000",
		16#022a# => X"00000000",
		16#022b# => X"00000000",
		16#022c# => X"00000000",
		16#022d# => X"00000000",
		16#022e# => X"00000000",
		16#022f# => X"00000000",
		16#0230# => X"00000000",
		16#0231# => X"00000000",
		16#0232# => X"00000000",
		16#0233# => X"00000000",
		16#0234# => X"00000000",
		16#0235# => X"00000000",
		16#0236# => X"00000000",
		16#0237# => X"00000000",
		16#0238# => X"00000000",
		16#0239# => X"00000000",
		16#023a# => X"00000000",
		16#023b# => X"00000000",
		16#023c# => X"00000000",
		16#023d# => X"00000000",
		16#023e# => X"00000000",
		16#023f# => X"00000000",
		16#0240# => X"00000000",
		16#0241# => X"00000000",
		16#0242# => X"00000000",
		16#0243# => X"00000000",
		16#0244# => X"00000000",
		16#0245# => X"00000000",
		16#0246# => X"00000000",
		16#0247# => X"00000000",
		16#0248# => X"00000000",
		16#0249# => X"00000000",
		16#024a# => X"00000000",
		16#024b# => X"00000000",
		16#024c# => X"00000000",
		16#024d# => X"00000000",
		16#024e# => X"00000000",
		16#024f# => X"00000000",
		16#0250# => X"00000000",
		16#0251# => X"00000000",
		16#0252# => X"00000000",
		16#0253# => X"00000000",
		16#0254# => X"00000000",
		16#0255# => X"00000000",
		16#0256# => X"00000000",
		16#0257# => X"00000000",
		16#0258# => X"00000000",
		16#0259# => X"00000000",
		16#025a# => X"00000000",
		16#025b# => X"00000000",
		16#025c# => X"00000000",
		16#025d# => X"00000000",
		16#025e# => X"00000000",
		16#025f# => X"00000000",
		16#0260# => X"00000000",
		16#0261# => X"00000000",
		16#0262# => X"00000000",
		16#0263# => X"00000000",
		16#0264# => X"00000000",
		16#0265# => X"00000000",
		16#0266# => X"00000000",
		16#0267# => X"00000000",
		16#0268# => X"00000000",
		16#0269# => X"00000000",
		16#026a# => X"00000000",
		16#026b# => X"00000000",
		16#026c# => X"00000000",
		16#026d# => X"00000000",
		16#026e# => X"00000000",
		16#026f# => X"00000000",
		16#0270# => X"00000000",
		16#0271# => X"00000000",
		16#0272# => X"00000000",
		16#0273# => X"00000000",
		16#0274# => X"00000000",
		16#0275# => X"00000000",
		16#0276# => X"00000000",
		16#0277# => X"00000000",
		16#0278# => X"00000000",
		16#0279# => X"00000000",
		16#027a# => X"00000000",
		16#027b# => X"00000000",
		16#027c# => X"00000000",
		16#027d# => X"00000000",
		16#027e# => X"00000000",
		16#027f# => X"00000000",
		16#0280# => X"00000000",
		16#0281# => X"00000000",
		16#0282# => X"00000000",
		16#0283# => X"00000000",
		16#0284# => X"00000000",
		16#0285# => X"00000000",
		16#0286# => X"00000000",
		16#0287# => X"00000000",
		16#0288# => X"00000000",
		16#0289# => X"00000000",
		16#028a# => X"00000000",
		16#028b# => X"00000000",
		16#028c# => X"00000000",
		16#028d# => X"00000000",
		16#028e# => X"00000000",
		16#028f# => X"00000000",
		16#0290# => X"00000000",
		16#0291# => X"00000000",
		16#0292# => X"00000000",
		16#0293# => X"00000000",
		16#0294# => X"00000000",
		16#0295# => X"00000000",
		16#0296# => X"00000000",
		16#0297# => X"00000000",
		16#0298# => X"00000000",
		16#0299# => X"00000000",
		16#029a# => X"00000000",
		16#029b# => X"00000000",
		16#029c# => X"00000000",
		16#029d# => X"00000000",
		16#029e# => X"00000000",
		16#029f# => X"00000000",
		16#02a0# => X"00000000",
		16#02a1# => X"00000000",
		16#02a2# => X"00000000",
		16#02a3# => X"00000000",
		16#02a4# => X"00000000",
		16#02a5# => X"00000000",
		16#02a6# => X"00000000",
		16#02a7# => X"00000000",
		16#02a8# => X"00000000",
		16#02a9# => X"00000000",
		16#02aa# => X"00000000",
		16#02ab# => X"00000000",
		16#02ac# => X"00000000",
		16#02ad# => X"00000000",
		16#02ae# => X"00000000",
		16#02af# => X"00000000",
		16#02b0# => X"00000000",
		16#02b1# => X"00000000",
		16#02b2# => X"00000000",
		16#02b3# => X"00000000",
		16#02b4# => X"00000000",
		16#02b5# => X"00000000",
		16#02b6# => X"00000000",
		16#02b7# => X"00000000",
		16#02b8# => X"00000000",
		16#02b9# => X"00000000",
		16#02ba# => X"00000000",
		16#02bb# => X"00000000",
		16#02bc# => X"00000000",
		16#02bd# => X"00000000",
		16#02be# => X"00000000",
		16#02bf# => X"00000000",
		16#02c0# => X"00000000",
		16#02c1# => X"00000000",
		16#02c2# => X"00000000",
		16#02c3# => X"00000000",
		16#02c4# => X"00000000",
		16#02c5# => X"00000000",
		16#02c6# => X"00000000",
		16#02c7# => X"00000000",
		16#02c8# => X"00000000",
		16#02c9# => X"00000000",
		16#02ca# => X"00000000",
		16#02cb# => X"00000000",
		16#02cc# => X"00000000",
		16#02cd# => X"00000000",
		16#02ce# => X"00000000",
		16#02cf# => X"00000000",
		16#02d0# => X"00000000",
		16#02d1# => X"00000000",
		16#02d2# => X"00000000",
		16#02d3# => X"00000000",
		16#02d4# => X"00000000",
		16#02d5# => X"00000000",
		16#02d6# => X"00000000",
		16#02d7# => X"00000000",
		16#02d8# => X"00000000",
		16#02d9# => X"00000000",
		16#02da# => X"00000000",
		16#02db# => X"00000000",
		16#02dc# => X"00000000",
		16#02dd# => X"00000000",
		16#02de# => X"00000000",
		16#02df# => X"00000000",
		16#02e0# => X"00000000",
		16#02e1# => X"00000000",
		16#02e2# => X"00000000",
		16#02e3# => X"00000000",
		16#02e4# => X"00000000",
		16#02e5# => X"00000000",
		16#02e6# => X"00000000",
		16#02e7# => X"00000000",
		16#02e8# => X"00000000",
		16#02e9# => X"00000000",
		16#02ea# => X"00000000",
		16#02eb# => X"00000000",
		16#02ec# => X"00000000",
		16#02ed# => X"00000000",
		16#02ee# => X"00000000",
		16#02ef# => X"00000000",
		16#02f0# => X"00000000",
		16#02f1# => X"00000000",
		16#02f2# => X"00000000",
		16#02f3# => X"00000000",
		16#02f4# => X"00000000",
		16#02f5# => X"00000000",
		16#02f6# => X"00000000",
		16#02f7# => X"00000000",
		16#02f8# => X"00000000",
		16#02f9# => X"00000000",
		16#02fa# => X"00000000",
		16#02fb# => X"00000000",
		16#02fc# => X"00000000",
		16#02fd# => X"00000000",
		16#02fe# => X"00000000",
		16#02ff# => X"00000000",
		16#0300# => X"24000000",
		16#0301# => X"00000000",
		16#0302# => X"00000000",
		16#0303# => X"00000000",
		16#0304# => X"00000000",
		16#0305# => X"00000000",
		16#0306# => X"00000000",
		16#0307# => X"00000000",
		16#0308# => X"00000000",
		16#0309# => X"00000000",
		16#030a# => X"00000000",
		16#030b# => X"00000000",
		16#030c# => X"00000000",
		16#030d# => X"00000000",
		16#030e# => X"00000000",
		16#030f# => X"00000000",
		16#0310# => X"00000000",
		16#0311# => X"00000000",
		16#0312# => X"00000000",
		16#0313# => X"00000000",
		16#0314# => X"00000000",
		16#0315# => X"00000000",
		16#0316# => X"00000000",
		16#0317# => X"00000000",
		16#0318# => X"00000000",
		16#0319# => X"00000000",
		16#031a# => X"00000000",
		16#031b# => X"00000000",
		16#031c# => X"00000000",
		16#031d# => X"00000000",
		16#031e# => X"00000000",
		16#031f# => X"00000000",
		16#0320# => X"00000000",
		16#0321# => X"00000000",
		16#0322# => X"00000000",
		16#0323# => X"00000000",
		16#0324# => X"00000000",
		16#0325# => X"00000000",
		16#0326# => X"00000000",
		16#0327# => X"00000000",
		16#0328# => X"00000000",
		16#0329# => X"00000000",
		16#032a# => X"00000000",
		16#032b# => X"00000000",
		16#032c# => X"00000000",
		16#032d# => X"00000000",
		16#032e# => X"00000000",
		16#032f# => X"00000000",
		16#0330# => X"00000000",
		16#0331# => X"00000000",
		16#0332# => X"00000000",
		16#0333# => X"00000000",
		16#0334# => X"00000000",
		16#0335# => X"00000000",
		16#0336# => X"00000000",
		16#0337# => X"00000000",
		16#0338# => X"00000000",
		16#0339# => X"00000000",
		16#033a# => X"00000000",
		16#033b# => X"00000000",
		16#033c# => X"00000000",
		16#033d# => X"00000000",
		16#033e# => X"00000000",
		16#033f# => X"00000000",
		16#0340# => X"00000000",
		16#0341# => X"00000000",
		16#0342# => X"00000000",
		16#0343# => X"00000000",
		16#0344# => X"00000000",
		16#0345# => X"00000000",
		16#0346# => X"00000000",
		16#0347# => X"00000000",
		16#0348# => X"00000000",
		16#0349# => X"00000000",
		16#034a# => X"00000000",
		16#034b# => X"00000000",
		16#034c# => X"00000000",
		16#034d# => X"00000000",
		16#034e# => X"00000000",
		16#034f# => X"00000000",
		16#0350# => X"00000000",
		16#0351# => X"00000000",
		16#0352# => X"00000000",
		16#0353# => X"00000000",
		16#0354# => X"00000000",
		16#0355# => X"00000000",
		16#0356# => X"00000000",
		16#0357# => X"00000000",
		16#0358# => X"00000000",
		16#0359# => X"00000000",
		16#035a# => X"00000000",
		16#035b# => X"00000000",
		16#035c# => X"00000000",
		16#035d# => X"00000000",
		16#035e# => X"00000000",
		16#035f# => X"00000000",
		16#0360# => X"00000000",
		16#0361# => X"00000000",
		16#0362# => X"00000000",
		16#0363# => X"00000000",
		16#0364# => X"00000000",
		16#0365# => X"00000000",
		16#0366# => X"00000000",
		16#0367# => X"00000000",
		16#0368# => X"00000000",
		16#0369# => X"00000000",
		16#036a# => X"00000000",
		16#036b# => X"00000000",
		16#036c# => X"00000000",
		16#036d# => X"00000000",
		16#036e# => X"00000000",
		16#036f# => X"00000000",
		16#0370# => X"00000000",
		16#0371# => X"00000000",
		16#0372# => X"00000000",
		16#0373# => X"00000000",
		16#0374# => X"00000000",
		16#0375# => X"00000000",
		16#0376# => X"00000000",
		16#0377# => X"00000000",
		16#0378# => X"00000000",
		16#0379# => X"00000000",
		16#037a# => X"00000000",
		16#037b# => X"00000000",
		16#037c# => X"00000000",
		16#037d# => X"00000000",
		16#037e# => X"00000000",
		16#037f# => X"00000000",
		16#0380# => X"18201500",
		16#0381# => X"d480081c",
		16#0382# => X"24000000",
		16#0383# => X"00000000",
		16#0384# => X"00000000",
		16#0385# => X"00000000",
		16#0386# => X"00000000",
		16#0387# => X"00000000",
		16#0388# => X"00000000",
		16#0389# => X"00000000",
		16#038a# => X"00000000",
		16#038b# => X"00000000",
		16#038c# => X"00000000",
		16#038d# => X"00000000",
		16#038e# => X"00000000",
		16#038f# => X"00000000",
		16#0390# => X"00000000",
		16#0391# => X"00000000",
		16#0392# => X"00000000",
		16#0393# => X"00000000",
		16#0394# => X"00000000",
		16#0395# => X"00000000",
		16#0396# => X"00000000",
		16#0397# => X"00000000",
		16#0398# => X"00000000",
		16#0399# => X"00000000",
		16#039a# => X"00000000",
		16#039b# => X"00000000",
		16#039c# => X"00000000",
		16#039d# => X"00000000",
		16#039e# => X"00000000",
		16#039f# => X"00000000",
		16#03a0# => X"00000000",
		16#03a1# => X"00000000",
		16#03a2# => X"00000000",
		16#03a3# => X"00000000",
		16#03a4# => X"00000000",
		16#03a5# => X"00000000",
		16#03a6# => X"00000000",
		16#03a7# => X"00000000",
		16#03a8# => X"00000000",
		16#03a9# => X"00000000",
		16#03aa# => X"00000000",
		16#03ab# => X"00000000",
		16#03ac# => X"00000000",
		16#03ad# => X"00000000",
		16#03ae# => X"00000000",
		16#03af# => X"00000000",
		16#03b0# => X"00000000",
		16#03b1# => X"00000000",
		16#03b2# => X"00000000",
		16#03b3# => X"00000000",
		16#03b4# => X"00000000",
		16#03b5# => X"00000000",
		16#03b6# => X"00000000",
		16#03b7# => X"00000000",
		16#03b8# => X"00000000",
		16#03b9# => X"00000000",
		16#03ba# => X"00000000",
		16#03bb# => X"00000000",
		16#03bc# => X"00000000",
		16#03bd# => X"00000000",
		16#03be# => X"00000000",
		16#03bf# => X"00000000",
		16#03c0# => X"00000000",
		16#03c1# => X"00000000",
		16#03c2# => X"00000000",
		16#03c3# => X"00000000",
		16#03c4# => X"00000000",
		16#03c5# => X"00000000",
		16#03c6# => X"00000000",
		16#03c7# => X"00000000",
		16#03c8# => X"00000000",
		16#03c9# => X"00000000",
		16#03ca# => X"00000000",
		16#03cb# => X"00000000",
		16#03cc# => X"00000000",
		16#03cd# => X"00000000",
		16#03ce# => X"00000000",
		16#03cf# => X"00000000",
		16#03d0# => X"00000000",
		16#03d1# => X"00000000",
		16#03d2# => X"00000000",
		16#03d3# => X"00000000",
		16#03d4# => X"00000000",
		16#03d5# => X"00000000",
		16#03d6# => X"00000000",
		16#03d7# => X"00000000",
		16#03d8# => X"00000000",
		16#03d9# => X"00000000",
		16#03da# => X"00000000",
		16#03db# => X"00000000",
		16#03dc# => X"00000000",
		16#03dd# => X"00000000",
		16#03de# => X"00000000",
		16#03df# => X"00000000",
		16#03e0# => X"00000000",
		16#03e1# => X"00000000",
		16#03e2# => X"00000000",
		16#03e3# => X"00000000",
		16#03e4# => X"00000000",
		16#03e5# => X"00000000",
		16#03e6# => X"00000000",
		16#03e7# => X"00000000",
		16#03e8# => X"00000000",
		16#03e9# => X"00000000",
		16#03ea# => X"00000000",
		16#03eb# => X"00000000",
		16#03ec# => X"00000000",
		16#03ed# => X"00000000",
		16#03ee# => X"00000000",
		16#03ef# => X"00000000",
		16#03f0# => X"00000000",
		16#03f1# => X"00000000",
		16#03f2# => X"00000000",
		16#03f3# => X"00000000",
		16#03f4# => X"00000000",
		16#03f5# => X"00000000",
		16#03f6# => X"00000000",
		16#03f7# => X"00000000",
		16#03f8# => X"00000000",
		16#03f9# => X"00000000",
		16#03fa# => X"00000000",
		16#03fb# => X"00000000",
		16#03fc# => X"00000000",
		16#03fd# => X"00000000",
		16#03fe# => X"00000000",
		16#03ff# => X"00000000",
		16#0400# => X"00000000",
		16#0401# => X"00000000",
		16#0402# => X"00000000",
		16#0403# => X"00000000",
		16#0404# => X"00000000",
		16#0405# => X"00000000",
		16#0406# => X"00000000",
		16#0407# => X"00000000",
		16#0408# => X"00000000",
		16#0409# => X"00000000",
		16#040a# => X"00000000",
		16#040b# => X"00000000",
		16#040c# => X"00000000",
		16#040d# => X"00000000",
		16#040e# => X"00000000",
		16#040f# => X"00000000",
		16#0410# => X"00000000",
		16#0411# => X"00000000",
		16#0412# => X"00000000",
		16#0413# => X"00000000",
		16#0414# => X"00000000",
		16#0415# => X"00000000",
		16#0416# => X"00000000",
		16#0417# => X"00000000",
		16#0418# => X"00000000",
		16#0419# => X"00000000",
		16#041a# => X"00000000",
		16#041b# => X"00000000",
		16#041c# => X"00000000",
		16#041d# => X"00000000",
		16#041e# => X"00000000",
		16#041f# => X"00000000",
		16#0420# => X"00000000",
		16#0421# => X"00000000",
		16#0422# => X"00000000",
		16#0423# => X"00000000",
		16#0424# => X"00000000",
		16#0425# => X"00000000",
		16#0426# => X"00000000",
		16#0427# => X"00000000",
		16#0428# => X"00000000",
		16#0429# => X"00000000",
		16#042a# => X"00000000",
		16#042b# => X"00000000",
		16#042c# => X"00000000",
		16#042d# => X"00000000",
		16#042e# => X"00000000",
		16#042f# => X"00000000",
		16#0430# => X"00000000",
		16#0431# => X"00000000",
		16#0432# => X"00000000",
		16#0433# => X"00000000",
		16#0434# => X"00000000",
		16#0435# => X"00000000",
		16#0436# => X"00000000",
		16#0437# => X"00000000",
		16#0438# => X"00000000",
		16#0439# => X"00000000",
		16#043a# => X"00000000",
		16#043b# => X"00000000",
		16#043c# => X"00000000",
		16#043d# => X"00000000",
		16#043e# => X"00000000",
		16#043f# => X"00000000",
		16#0440# => X"00000000",
		16#0441# => X"00000000",
		16#0442# => X"00000000",
		16#0443# => X"00000000",
		16#0444# => X"00000000",
		16#0445# => X"00000000",
		16#0446# => X"00000000",
		16#0447# => X"00000000",
		16#0448# => X"00000000",
		16#0449# => X"00000000",
		16#044a# => X"00000000",
		16#044b# => X"00000000",
		16#044c# => X"00000000",
		16#044d# => X"00000000",
		16#044e# => X"00000000",
		16#044f# => X"00000000",
		16#0450# => X"00000000",
		16#0451# => X"00000000",
		16#0452# => X"00000000",
		16#0453# => X"00000000",
		16#0454# => X"00000000",
		16#0455# => X"00000000",
		16#0456# => X"00000000",
		16#0457# => X"00000000",
		16#0458# => X"00000000",
		16#0459# => X"00000000",
		16#045a# => X"00000000",
		16#045b# => X"00000000",
		16#045c# => X"00000000",
		16#045d# => X"00000000",
		16#045e# => X"00000000",
		16#045f# => X"00000000",
		16#0460# => X"00000000",
		16#0461# => X"00000000",
		16#0462# => X"00000000",
		16#0463# => X"00000000",
		16#0464# => X"00000000",
		16#0465# => X"00000000",
		16#0466# => X"00000000",
		16#0467# => X"00000000",
		16#0468# => X"00000000",
		16#0469# => X"00000000",
		16#046a# => X"00000000",
		16#046b# => X"00000000",
		16#046c# => X"00000000",
		16#046d# => X"00000000",
		16#046e# => X"00000000",
		16#046f# => X"00000000",
		16#0470# => X"00000000",
		16#0471# => X"00000000",
		16#0472# => X"00000000",
		16#0473# => X"00000000",
		16#0474# => X"00000000",
		16#0475# => X"00000000",
		16#0476# => X"00000000",
		16#0477# => X"00000000",
		16#0478# => X"00000000",
		16#0479# => X"00000000",
		16#047a# => X"00000000",
		16#047b# => X"00000000",
		16#047c# => X"00000000",
		16#047d# => X"00000000",
		16#047e# => X"00000000",
		16#047f# => X"00000000",
		16#0480# => X"00000000",
		16#0481# => X"00000000",
		16#0482# => X"00000000",
		16#0483# => X"00000000",
		16#0484# => X"00000000",
		16#0485# => X"00000000",
		16#0486# => X"00000000",
		16#0487# => X"00000000",
		16#0488# => X"00000000",
		16#0489# => X"00000000",
		16#048a# => X"00000000",
		16#048b# => X"00000000",
		16#048c# => X"00000000",
		16#048d# => X"00000000",
		16#048e# => X"00000000",
		16#048f# => X"00000000",
		16#0490# => X"00000000",
		16#0491# => X"00000000",
		16#0492# => X"00000000",
		16#0493# => X"00000000",
		16#0494# => X"00000000",
		16#0495# => X"00000000",
		16#0496# => X"00000000",
		16#0497# => X"00000000",
		16#0498# => X"00000000",
		16#0499# => X"00000000",
		16#049a# => X"00000000",
		16#049b# => X"00000000",
		16#049c# => X"00000000",
		16#049d# => X"00000000",
		16#049e# => X"00000000",
		16#049f# => X"00000000",
		16#04a0# => X"00000000",
		16#04a1# => X"00000000",
		16#04a2# => X"00000000",
		16#04a3# => X"00000000",
		16#04a4# => X"00000000",
		16#04a5# => X"00000000",
		16#04a6# => X"00000000",
		16#04a7# => X"00000000",
		16#04a8# => X"00000000",
		16#04a9# => X"00000000",
		16#04aa# => X"00000000",
		16#04ab# => X"00000000",
		16#04ac# => X"00000000",
		16#04ad# => X"00000000",
		16#04ae# => X"00000000",
		16#04af# => X"00000000",
		16#04b0# => X"00000000",
		16#04b1# => X"00000000",
		16#04b2# => X"00000000",
		16#04b3# => X"00000000",
		16#04b4# => X"00000000",
		16#04b5# => X"00000000",
		16#04b6# => X"00000000",
		16#04b7# => X"00000000",
		16#04b8# => X"00000000",
		16#04b9# => X"00000000",
		16#04ba# => X"00000000",
		16#04bb# => X"00000000",
		16#04bc# => X"00000000",
		16#04bd# => X"00000000",
		16#04be# => X"00000000",
		16#04bf# => X"00000000",
		16#04c0# => X"00000000",
		16#04c1# => X"00000000",
		16#04c2# => X"00000000",
		16#04c3# => X"00000000",
		16#04c4# => X"00000000",
		16#04c5# => X"00000000",
		16#04c6# => X"00000000",
		16#04c7# => X"00000000",
		16#04c8# => X"00000000",
		16#04c9# => X"00000000",
		16#04ca# => X"00000000",
		16#04cb# => X"00000000",
		16#04cc# => X"00000000",
		16#04cd# => X"00000000",
		16#04ce# => X"00000000",
		16#04cf# => X"00000000",
		16#04d0# => X"00000000",
		16#04d1# => X"00000000",
		16#04d2# => X"00000000",
		16#04d3# => X"00000000",
		16#04d4# => X"00000000",
		16#04d5# => X"00000000",
		16#04d6# => X"00000000",
		16#04d7# => X"00000000",
		16#04d8# => X"00000000",
		16#04d9# => X"00000000",
		16#04da# => X"00000000",
		16#04db# => X"00000000",
		16#04dc# => X"00000000",
		16#04dd# => X"00000000",
		16#04de# => X"00000000",
		16#04df# => X"00000000",
		16#04e0# => X"00000000",
		16#04e1# => X"00000000",
		16#04e2# => X"00000000",
		16#04e3# => X"00000000",
		16#04e4# => X"00000000",
		16#04e5# => X"00000000",
		16#04e6# => X"00000000",
		16#04e7# => X"00000000",
		16#04e8# => X"00000000",
		16#04e9# => X"00000000",
		16#04ea# => X"00000000",
		16#04eb# => X"00000000",
		16#04ec# => X"00000000",
		16#04ed# => X"00000000",
		16#04ee# => X"00000000",
		16#04ef# => X"00000000",
		16#04f0# => X"00000000",
		16#04f1# => X"00000000",
		16#04f2# => X"00000000",
		16#04f3# => X"00000000",
		16#04f4# => X"00000000",
		16#04f5# => X"00000000",
		16#04f6# => X"00000000",
		16#04f7# => X"00000000",
		16#04f8# => X"00000000",
		16#04f9# => X"00000000",
		16#04fa# => X"00000000",
		16#04fb# => X"00000000",
		16#04fc# => X"00000000",
		16#04fd# => X"00000000",
		16#04fe# => X"00000000",
		16#04ff# => X"00000000",
		16#0500# => X"00000000",
		16#0501# => X"00000000",
		16#0502# => X"00000000",
		16#0503# => X"00000000",
		16#0504# => X"00000000",
		16#0505# => X"00000000",
		16#0506# => X"00000000",
		16#0507# => X"00000000",
		16#0508# => X"00000000",
		16#0509# => X"00000000",
		16#050a# => X"00000000",
		16#050b# => X"00000000",
		16#050c# => X"00000000",
		16#050d# => X"00000000",
		16#050e# => X"00000000",
		16#050f# => X"00000000",
		16#0510# => X"00000000",
		16#0511# => X"00000000",
		16#0512# => X"00000000",
		16#0513# => X"00000000",
		16#0514# => X"00000000",
		16#0515# => X"00000000",
		16#0516# => X"00000000",
		16#0517# => X"00000000",
		16#0518# => X"00000000",
		16#0519# => X"00000000",
		16#051a# => X"00000000",
		16#051b# => X"00000000",
		16#051c# => X"00000000",
		16#051d# => X"00000000",
		16#051e# => X"00000000",
		16#051f# => X"00000000",
		16#0520# => X"00000000",
		16#0521# => X"00000000",
		16#0522# => X"00000000",
		16#0523# => X"00000000",
		16#0524# => X"00000000",
		16#0525# => X"00000000",
		16#0526# => X"00000000",
		16#0527# => X"00000000",
		16#0528# => X"00000000",
		16#0529# => X"00000000",
		16#052a# => X"00000000",
		16#052b# => X"00000000",
		16#052c# => X"00000000",
		16#052d# => X"00000000",
		16#052e# => X"00000000",
		16#052f# => X"00000000",
		16#0530# => X"00000000",
		16#0531# => X"00000000",
		16#0532# => X"00000000",
		16#0533# => X"00000000",
		16#0534# => X"00000000",
		16#0535# => X"00000000",
		16#0536# => X"00000000",
		16#0537# => X"00000000",
		16#0538# => X"00000000",
		16#0539# => X"00000000",
		16#053a# => X"00000000",
		16#053b# => X"00000000",
		16#053c# => X"00000000",
		16#053d# => X"00000000",
		16#053e# => X"00000000",
		16#053f# => X"00000000",
		16#0540# => X"00000000",
		16#0541# => X"00000000",
		16#0542# => X"00000000",
		16#0543# => X"00000000",
		16#0544# => X"00000000",
		16#0545# => X"00000000",
		16#0546# => X"00000000",
		16#0547# => X"00000000",
		16#0548# => X"00000000",
		16#0549# => X"00000000",
		16#054a# => X"00000000",
		16#054b# => X"00000000",
		16#054c# => X"00000000",
		16#054d# => X"00000000",
		16#054e# => X"00000000",
		16#054f# => X"00000000",
		16#0550# => X"00000000",
		16#0551# => X"00000000",
		16#0552# => X"00000000",
		16#0553# => X"00000000",
		16#0554# => X"00000000",
		16#0555# => X"00000000",
		16#0556# => X"00000000",
		16#0557# => X"00000000",
		16#0558# => X"00000000",
		16#0559# => X"00000000",
		16#055a# => X"00000000",
		16#055b# => X"00000000",
		16#055c# => X"00000000",
		16#055d# => X"00000000",
		16#055e# => X"00000000",
		16#055f# => X"00000000",
		16#0560# => X"00000000",
		16#0561# => X"00000000",
		16#0562# => X"00000000",
		16#0563# => X"00000000",
		16#0564# => X"00000000",
		16#0565# => X"00000000",
		16#0566# => X"00000000",
		16#0567# => X"00000000",
		16#0568# => X"00000000",
		16#0569# => X"00000000",
		16#056a# => X"00000000",
		16#056b# => X"00000000",
		16#056c# => X"00000000",
		16#056d# => X"00000000",
		16#056e# => X"00000000",
		16#056f# => X"00000000",
		16#0570# => X"00000000",
		16#0571# => X"00000000",
		16#0572# => X"00000000",
		16#0573# => X"00000000",
		16#0574# => X"00000000",
		16#0575# => X"00000000",
		16#0576# => X"00000000",
		16#0577# => X"00000000",
		16#0578# => X"00000000",
		16#0579# => X"00000000",
		16#057a# => X"00000000",
		16#057b# => X"00000000",
		16#057c# => X"00000000",
		16#057d# => X"00000000",
		16#057e# => X"00000000",
		16#057f# => X"00000000",
		16#0580# => X"00000000",
		16#0581# => X"00000000",
		16#0582# => X"00000000",
		16#0583# => X"00000000",
		16#0584# => X"00000000",
		16#0585# => X"00000000",
		16#0586# => X"00000000",
		16#0587# => X"00000000",
		16#0588# => X"00000000",
		16#0589# => X"00000000",
		16#058a# => X"00000000",
		16#058b# => X"00000000",
		16#058c# => X"00000000",
		16#058d# => X"00000000",
		16#058e# => X"00000000",
		16#058f# => X"00000000",
		16#0590# => X"00000000",
		16#0591# => X"00000000",
		16#0592# => X"00000000",
		16#0593# => X"00000000",
		16#0594# => X"00000000",
		16#0595# => X"00000000",
		16#0596# => X"00000000",
		16#0597# => X"00000000",
		16#0598# => X"00000000",
		16#0599# => X"00000000",
		16#059a# => X"00000000",
		16#059b# => X"00000000",
		16#059c# => X"00000000",
		16#059d# => X"00000000",
		16#059e# => X"00000000",
		16#059f# => X"00000000",
		16#05a0# => X"00000000",
		16#05a1# => X"00000000",
		16#05a2# => X"00000000",
		16#05a3# => X"00000000",
		16#05a4# => X"00000000",
		16#05a5# => X"00000000",
		16#05a6# => X"00000000",
		16#05a7# => X"00000000",
		16#05a8# => X"00000000",
		16#05a9# => X"00000000",
		16#05aa# => X"00000000",
		16#05ab# => X"00000000",
		16#05ac# => X"00000000",
		16#05ad# => X"00000000",
		16#05ae# => X"00000000",
		16#05af# => X"00000000",
		16#05b0# => X"00000000",
		16#05b1# => X"00000000",
		16#05b2# => X"00000000",
		16#05b3# => X"00000000",
		16#05b4# => X"00000000",
		16#05b5# => X"00000000",
		16#05b6# => X"00000000",
		16#05b7# => X"00000000",
		16#05b8# => X"00000000",
		16#05b9# => X"00000000",
		16#05ba# => X"00000000",
		16#05bb# => X"00000000",
		16#05bc# => X"00000000",
		16#05bd# => X"00000000",
		16#05be# => X"00000000",
		16#05bf# => X"00000000",
		16#05c0# => X"ffffffff",
		16#05c1# => X"ffffffff",
		16#05c2# => X"ffffffff",
		16#05c3# => X"ffffffff",
		16#05c4# => X"ffffffff",
		16#05c5# => X"ffffffff",
		16#05c6# => X"ffffffff",
		16#05c7# => X"ffffffff",
		16#05c8# => X"ffffffff",
		16#05c9# => X"ffffffff",
		16#05ca# => X"deadbeef",
		16#05cb# => X"00000000",
		16#05cc# => X"00000000",
		16#05cd# => X"00000000",
		16#05ce# => X"00000000",
		16#05cf# => X"00000000",
		16#05d0# => X"00000000",
		16#05d1# => X"00000000",
		16#05d2# => X"00000000",
		16#05d3# => X"00000000",
		16#05d4# => X"00000000",
		16#05d5# => X"00000000",
		16#05d6# => X"00000000",
		16#05d7# => X"00000000",
		16#05d8# => X"00000000",
		16#05d9# => X"00000000",
		16#05da# => X"00000000",
		16#05db# => X"00000000",
		16#05dc# => X"00000000",
		16#05dd# => X"00000000",
		16#05de# => X"00000000",
		16#05df# => X"00000000",
		16#05e0# => X"00000000",
		16#05e1# => X"00000000",
		16#05e2# => X"00000000",
		16#05e3# => X"00000000",
		16#05e4# => X"00000000",
		16#05e5# => X"00000000",
		16#05e6# => X"00000000",
		16#05e7# => X"00000000",
		16#05e8# => X"00000000",
		16#05e9# => X"00000000",
		16#05ea# => X"00000000",
		16#05eb# => X"00000000",
		16#05ec# => X"00000000",
		16#05ed# => X"00000000",
		16#05ee# => X"00000000",
		16#05ef# => X"00000000",
		16#05f0# => X"00000000",
		16#05f1# => X"00000000",
		16#05f2# => X"00000000",
		16#05f3# => X"00000000",
		16#05f4# => X"00000000",
		16#05f5# => X"00000000",
		16#05f6# => X"00000000",
		16#05f7# => X"00000000",
		16#05f8# => X"00000000",
		16#05f9# => X"00000000",
		16#05fa# => X"00000000",
		16#05fb# => X"00000000",
		16#05fc# => X"00000000",
		16#05fd# => X"00000000",
		16#05fe# => X"00000000",
		16#05ff# => X"00000000",
		16#0600# => X"00000000",
		16#0601# => X"00000000",
		16#0602# => X"00000000",
		16#0603# => X"00000000",
		16#0604# => X"00000000",
		16#0605# => X"00000000",
		16#0606# => X"00000000",
		16#0607# => X"00000000",
		16#0608# => X"00000000",
		16#0609# => X"00000000",
		16#060a# => X"00000000",
		16#060b# => X"00000000",
		16#060c# => X"00000000",
		16#060d# => X"00000000",
		16#060e# => X"00000000",
		16#060f# => X"00000000",
		16#0610# => X"00000000",
		16#0611# => X"00000000",
		16#0612# => X"00000000",
		16#0613# => X"00000000",
		16#0614# => X"00000000",
		16#0615# => X"00000000",
		16#0616# => X"00000000",
		16#0617# => X"00000000",
		16#0618# => X"00000000",
		16#0619# => X"00000000",
		16#061a# => X"00000000",
		16#061b# => X"00000000",
		16#061c# => X"00000000",
		16#061d# => X"00000000",
		16#061e# => X"00000000",
		16#061f# => X"00000000",
		16#0620# => X"00000000",
		16#0621# => X"00000000",
		16#0622# => X"00000000",
		16#0623# => X"00000000",
		16#0624# => X"00000000",
		16#0625# => X"00000000",
		16#0626# => X"00000000",
		16#0627# => X"00000000",
		16#0628# => X"00000000",
		16#0629# => X"00000000",
		16#062a# => X"00000000",
		16#062b# => X"00000000",
		16#062c# => X"00000000",
		16#062d# => X"00000000",
		16#062e# => X"00000000",
		16#062f# => X"00000000",
		16#0630# => X"00000000",
		16#0631# => X"00000000",
		16#0632# => X"00000000",
		16#0633# => X"00000000",
		16#0634# => X"00000000",
		16#0635# => X"00000000",
		16#0636# => X"00000000",
		16#0637# => X"00000000",
		16#0638# => X"00000000",
		16#0639# => X"00000000",
		16#063a# => X"00000000",
		16#063b# => X"00000000",
		16#063c# => X"00000000",
		16#063d# => X"00000000",
		16#063e# => X"00000000",
		16#063f# => X"00000000",
		16#0640# => X"00000000",
		16#0641# => X"00000000",
		16#0642# => X"00000000",
		16#0643# => X"00000000",
		16#0644# => X"00000000",
		16#0645# => X"00000000",
		16#0646# => X"00000000",
		16#0647# => X"00000000",
		16#0648# => X"00000000",
		16#0649# => X"00000000",
		16#064a# => X"00000000",
		16#064b# => X"00000000",
		16#064c# => X"00000000",
		16#064d# => X"00000000",
		16#064e# => X"00000000",
		16#064f# => X"00000000",
		16#0650# => X"00000000",
		16#0651# => X"00000000",
		16#0652# => X"00000000",
		16#0653# => X"00000000",
		16#0654# => X"00000000",
		16#0655# => X"00000000",
		16#0656# => X"00000000",
		16#0657# => X"00000000",
		16#0658# => X"00000000",
		16#0659# => X"00000000",
		16#065a# => X"00000000",
		16#065b# => X"00000000",
		16#065c# => X"00000000",
		16#065d# => X"00000000",
		16#065e# => X"00000000",
		16#065f# => X"00000000",
		16#0660# => X"00000000",
		16#0661# => X"00000000",
		16#0662# => X"00000000",
		16#0663# => X"00000000",
		16#0664# => X"00000000",
		16#0665# => X"00000000",
		16#0666# => X"00000000",
		16#0667# => X"00000000",
		16#0668# => X"00000000",
		16#0669# => X"00000000",
		16#066a# => X"00000000",
		16#066b# => X"00000000",
		16#066c# => X"00000000",
		16#066d# => X"00000000",
		16#066e# => X"00000000",
		16#066f# => X"00000000",
		16#0670# => X"00000000",
		16#0671# => X"00000000",
		16#0672# => X"00000000",
		16#0673# => X"00000000",
		16#0674# => X"00000000",
		16#0675# => X"00000000",
		16#0676# => X"00000000",
		16#0677# => X"00000000",
		16#0678# => X"00000000",
		16#0679# => X"00000000",
		16#067a# => X"00000000",
		16#067b# => X"00000000",
		16#067c# => X"00000000",
		16#067d# => X"00000000",
		16#067e# => X"00000000",
		16#067f# => X"00000000",
		16#0680# => X"00000000",
		16#0681# => X"00000000",
		16#0682# => X"00000000",
		16#0683# => X"00000000",
		16#0684# => X"00000000",
		16#0685# => X"00000000",
		16#0686# => X"00000000",
		16#0687# => X"00000000",
		16#0688# => X"00000000",
		16#0689# => X"00000000",
		16#068a# => X"00000000",
		16#068b# => X"00000000",
		16#068c# => X"00000000",
		16#068d# => X"00000000",
		16#068e# => X"00000000",
		16#068f# => X"00000000",
		16#0690# => X"00000000",
		16#0691# => X"00000000",
		16#0692# => X"00000000",
		16#0693# => X"00000000",
		16#0694# => X"00000000",
		16#0695# => X"00000000",
		16#0696# => X"00000000",
		16#0697# => X"00000000",
		16#0698# => X"00000000",
		16#0699# => X"00000000",
		16#069a# => X"00000000",
		16#069b# => X"00000000",
		16#069c# => X"00000000",
		16#069d# => X"00000000",
		16#069e# => X"00000000",
		16#069f# => X"00000000",
		16#06a0# => X"00000000",
		16#06a1# => X"00000000",
		16#06a2# => X"00000000",
		16#06a3# => X"00000000",
		16#06a4# => X"00000000",
		16#06a5# => X"00000000",
		16#06a6# => X"00000000",
		16#06a7# => X"00000000",
		16#06a8# => X"00000000",
		16#06a9# => X"00000000",
		16#06aa# => X"00000000",
		16#06ab# => X"00000000",
		16#06ac# => X"00000000",
		16#06ad# => X"00000000",
		16#06ae# => X"00000000",
		16#06af# => X"00000000",
		16#06b0# => X"00000000",
		16#06b1# => X"00000000",
		16#06b2# => X"00000000",
		16#06b3# => X"00000000",
		16#06b4# => X"00000000",
		16#06b5# => X"00000000",
		16#06b6# => X"00000000",
		16#06b7# => X"00000000",
		16#06b8# => X"00000000",
		16#06b9# => X"00000000",
		16#06ba# => X"00000000",
		16#06bb# => X"00000000",
		16#06bc# => X"00000000",
		16#06bd# => X"00000000",
		16#06be# => X"00000000",
		16#06bf# => X"00000000",
		16#06c0# => X"00000000",
		16#06c1# => X"00000000",
		16#06c2# => X"00000000",
		16#06c3# => X"00000000",
		16#06c4# => X"00000000",
		16#06c5# => X"00000000",
		16#06c6# => X"00000000",
		16#06c7# => X"00000000",
		16#06c8# => X"00000000",
		16#06c9# => X"00000000",
		16#06ca# => X"00000000",
		16#06cb# => X"00000000",
		16#06cc# => X"00000000",
		16#06cd# => X"00000000",
		16#06ce# => X"00000000",
		16#06cf# => X"00000000",
		16#06d0# => X"00000000",
		16#06d1# => X"00000000",
		16#06d2# => X"00000000",
		16#06d3# => X"00000000",
		16#06d4# => X"00000000",
		16#06d5# => X"00000000",
		16#06d6# => X"00000000",
		16#06d7# => X"00000000",
		16#06d8# => X"00000000",
		16#06d9# => X"00000000",
		16#06da# => X"00000000",
		16#06db# => X"00000000",
		16#06dc# => X"00000000",
		16#06dd# => X"00000000",
		16#06de# => X"00000000",
		16#06df# => X"00000000",
		16#06e0# => X"00000000",
		16#06e1# => X"00000000",
		16#06e2# => X"00000000",
		16#06e3# => X"00000000",
		16#06e4# => X"00000000",
		16#06e5# => X"00000000",
		16#06e6# => X"00000000",
		16#06e7# => X"00000000",
		16#06e8# => X"00000000",
		16#06e9# => X"00000000",
		16#06ea# => X"00000000",
		16#06eb# => X"00000000",
		16#06ec# => X"00000000",
		16#06ed# => X"00000000",
		16#06ee# => X"00000000",
		16#06ef# => X"00000000",
		16#06f0# => X"00000000",
		16#06f1# => X"00000000",
		16#06f2# => X"00000000",
		16#06f3# => X"00000000",
		16#06f4# => X"00000000",
		16#06f5# => X"00000000",
		16#06f6# => X"00000000",
		16#06f7# => X"00000000",
		16#06f8# => X"00000000",
		16#06f9# => X"00000000",
		16#06fa# => X"00000000",
		16#06fb# => X"00000000",
		16#06fc# => X"00000000",
		16#06fd# => X"00000000",
		16#06fe# => X"00000000",
		16#06ff# => X"00000000",
		16#0700# => X"00000000",
		16#0701# => X"00000000",
		16#0702# => X"00000000",
		16#0703# => X"00000000",
		16#0704# => X"00000000",
		16#0705# => X"00000000",
		16#0706# => X"00000000",
		16#0707# => X"00000000",
		16#0708# => X"00000000",
		16#0709# => X"00000000",
		16#070a# => X"00000000",
		16#070b# => X"00000000",
		16#070c# => X"00000000",
		16#070d# => X"00000000",
		16#070e# => X"00000000",
		16#070f# => X"00000000",
		16#0710# => X"00000000",
		16#0711# => X"00000000",
		16#0712# => X"00000000",
		16#0713# => X"00000000",
		16#0714# => X"00000000",
		16#0715# => X"00000000",
		16#0716# => X"00000000",
		16#0717# => X"00000000",
		16#0718# => X"00000000",
		16#0719# => X"00000000",
		16#071a# => X"00000000",
		16#071b# => X"00000000",
		16#071c# => X"00000000",
		16#071d# => X"00000000",
		16#071e# => X"00000000",
		16#071f# => X"00000000",
		16#0720# => X"00000000",
		16#0721# => X"00000000",
		16#0722# => X"00000000",
		16#0723# => X"00000000",
		16#0724# => X"00000000",
		16#0725# => X"00000000",
		16#0726# => X"00000000",
		16#0727# => X"00000000",
		16#0728# => X"00000000",
		16#0729# => X"00000000",
		16#072a# => X"00000000",
		16#072b# => X"00000000",
		16#072c# => X"00000000",
		16#072d# => X"00000000",
		16#072e# => X"00000000",
		16#072f# => X"00000000",
		16#0730# => X"00000000",
		16#0731# => X"00000000",
		16#0732# => X"00000000",
		16#0733# => X"00000000",
		16#0734# => X"00000000",
		16#0735# => X"00000000",
		16#0736# => X"00000000",
		16#0737# => X"00000000",
		16#0738# => X"00000000",
		16#0739# => X"00000000",
		16#073a# => X"00000000",
		16#073b# => X"00000000",
		16#073c# => X"00000000",
		16#073d# => X"00000000",
		16#073e# => X"00000000",
		16#073f# => X"00000000",
		16#0740# => X"00000000",
		16#0741# => X"00000000",
		16#0742# => X"00000000",
		16#0743# => X"00000000",
		16#0744# => X"00000000",
		16#0745# => X"00000000",
		16#0746# => X"00000000",
		16#0747# => X"00000000",
		16#0748# => X"00000000",
		16#0749# => X"00000000",
		16#074a# => X"00000000",
		16#074b# => X"00000000",
		16#074c# => X"00000000",
		16#074d# => X"00000000",
		16#074e# => X"00000000",
		16#074f# => X"00000000",
		16#0750# => X"00000000",
		16#0751# => X"00000000",
		16#0752# => X"00000000",
		16#0753# => X"00000000",
		16#0754# => X"00000000",
		16#0755# => X"00000000",
		16#0756# => X"00000000",
		16#0757# => X"00000000",
		16#0758# => X"00000000",
		16#0759# => X"00000000",
		16#075a# => X"00000000",
		16#075b# => X"00000000",
		16#075c# => X"00000000",
		16#075d# => X"00000000",
		16#075e# => X"00000000",
		16#075f# => X"00000000",
		16#0760# => X"00000000",
		16#0761# => X"00000000",
		16#0762# => X"00000000",
		16#0763# => X"00000000",
		16#0764# => X"00000000",
		16#0765# => X"00000000",
		16#0766# => X"00000000",
		16#0767# => X"00000000",
		16#0768# => X"00000000",
		16#0769# => X"00000000",
		16#076a# => X"00000000",
		16#076b# => X"00000000",
		16#076c# => X"00000000",
		16#076d# => X"00000000",
		16#076e# => X"00000000",
		16#076f# => X"00000000",
		16#0770# => X"00000000",
		16#0771# => X"00000000",
		16#0772# => X"00000000",
		16#0773# => X"00000000",
		16#0774# => X"00000000",
		16#0775# => X"00000000",
		16#0776# => X"00000000",
		16#0777# => X"00000000",
		16#0778# => X"00000000",
		16#0779# => X"00000000",
		16#077a# => X"00000000",
		16#077b# => X"00000000",
		16#077c# => X"00000000",
		16#077d# => X"00000000",
		16#077e# => X"00000000",
		16#077f# => X"00000000",
		16#0780# => X"00000000",
		16#0781# => X"00000000",
		16#0782# => X"00000000",
		16#0783# => X"00000000",
		16#0784# => X"00000000",
		16#0785# => X"00000000",
		16#0786# => X"00000000",
		16#0787# => X"00000000",
		16#0788# => X"00000000",
		16#0789# => X"00000000",
		16#078a# => X"00000000",
		16#078b# => X"00000000",
		16#078c# => X"00000000",
		16#078d# => X"00000000",
		16#078e# => X"00000000",
		16#078f# => X"00000000",
		16#0790# => X"00000000",
		16#0791# => X"00000000",
		16#0792# => X"00000000",
		16#0793# => X"00000000",
		16#0794# => X"00000000",
		16#0795# => X"00000000",
		16#0796# => X"00000000",
		16#0797# => X"00000000",
		16#0798# => X"00000000",
		16#0799# => X"00000000",
		16#079a# => X"00000000",
		16#079b# => X"00000000",
		16#079c# => X"00000000",
		16#079d# => X"00000000",
		16#079e# => X"00000000",
		16#079f# => X"00000000",
		16#07a0# => X"00000000",
		16#07a1# => X"00000000",
		16#07a2# => X"00000000",
		16#07a3# => X"00000000",
		16#07a4# => X"00000000",
		16#07a5# => X"00000000",
		16#07a6# => X"00000000",
		16#07a7# => X"00000000",
		16#07a8# => X"00000000",
		16#07a9# => X"00000000",
		16#07aa# => X"00000000",
		16#07ab# => X"00000000",
		16#07ac# => X"00000000",
		16#07ad# => X"00000000",
		16#07ae# => X"00000000",
		16#07af# => X"00000000",
		16#07b0# => X"00000000",
		16#07b1# => X"00000000",
		16#07b2# => X"00000000",
		16#07b3# => X"00000000",
		16#07b4# => X"00000000",
		16#07b5# => X"00000000",
		16#07b6# => X"00000000",
		16#07b7# => X"00000000",
		16#07b8# => X"00000000",
		16#07b9# => X"00000000",
		16#07ba# => X"00000000",
		16#07bb# => X"00000000",
		16#07bc# => X"00000000",
		16#07bd# => X"00000000",
		16#07be# => X"00000000",
		16#07bf# => X"00000000",
		16#07c0# => X"00000000",
		16#07c1# => X"00000000",
		16#07c2# => X"00000000",
		16#07c3# => X"00000000",
		16#07c4# => X"00000000",
		16#07c5# => X"00000000",
		16#07c6# => X"00000000",
		16#07c7# => X"00000000",
		16#07c8# => X"00000000",
		16#07c9# => X"00000000",
		16#07ca# => X"00000000",
		16#07cb# => X"00000000",
		16#07cc# => X"00000000",
		16#07cd# => X"00000000",
		16#07ce# => X"00000000",
		16#07cf# => X"00000000",
		16#07d0# => X"00000000",
		16#07d1# => X"00000000",
		16#07d2# => X"00000000",
		16#07d3# => X"00000000",
		16#07d4# => X"00000000",
		16#07d5# => X"00000000",
		16#07d6# => X"00000000",
		16#07d7# => X"00000000",
		16#07d8# => X"00000000",
		16#07d9# => X"00000000",
		16#07da# => X"00000000",
		16#07db# => X"00000000",
		16#07dc# => X"00000000",
		16#07dd# => X"00000000",
		16#07de# => X"00000000",
		16#07df# => X"00000000",
		16#07e0# => X"00000000",
		16#07e1# => X"00000000",
		16#07e2# => X"00000000",
		16#07e3# => X"00000000",
		16#07e4# => X"00000000",
		16#07e5# => X"00000000",
		16#07e6# => X"00000000",
		16#07e7# => X"00000000",
		16#07e8# => X"00000000",
		16#07e9# => X"00000000",
		16#07ea# => X"00000000",
		16#07eb# => X"00000000",
		16#07ec# => X"00000000",
		16#07ed# => X"00000000",
		16#07ee# => X"00000000",
		16#07ef# => X"00000000",
		16#07f0# => X"00000000",
		16#07f1# => X"00000000",
		16#07f2# => X"00000000",
		16#07f3# => X"00000000",
		16#07f4# => X"00000000",
		16#07f5# => X"00000000",
		16#07f6# => X"00000000",
		16#07f7# => X"00000000",
		16#07f8# => X"00000000",
		16#07f9# => X"00000000",
		16#07fa# => X"00000000",
		16#07fb# => X"00000000",
		16#07fc# => X"00000000",
		16#07fd# => X"00000000",
		16#07fe# => X"00000000",
		16#07ff# => X"00000000",
		16#0800# => X"15000000",
		16#0801# => X"18200000",
		16#0802# => X"a8208005",
		16#0803# => X"c0000811",
		16#0804# => X"20000000",
		16#0805# => X"9c000000",
		16#0806# => X"15000000",
		16#0807# => X"21000000",
		16#0808# => X"15000000",
		16#0809# => X"d4000001",
		16#080a# => X"15000000",
		16#080b# => X"c8000014",
		16#080c# => X"15000000",
		16#080d# => X"00000001",
		16#080e# => X"1840cafe",
		16#080f# => X"a842babe",
		16#0810# => X"d4401700",
		16#0811# => X"18200000",
		16#0812# => X"a8211700",
		16#0813# => X"84210000",
		16#0814# => X"e0611005",
		16#0815# => X"98801700",
		16#0816# => X"1840ffff",
		16#0817# => X"a842cafe",
		16#0818# => X"e0a41005",
		16#0819# => X"e0632804",
		16#081a# => X"94a01702",
		16#081b# => X"18400000",
		16#081c# => X"a842babe",
		16#081d# => X"e0a51005",
		16#081e# => X"e0632804",
		16#081f# => X"18200000",
		16#0820# => X"a8211700",
		16#0821# => X"90c10000",
		16#0822# => X"90e10002",
		16#0823# => X"91010003",
		16#0824# => X"8d210001",
		16#0825# => X"8d410002",
		16#0826# => X"8d610003",
		16#0827# => X"e1864805",
		16#0828# => X"e1a75805",
		16#0829# => X"e1c85005",
		16#082a# => X"19e0ffff",
		16#082b# => X"a9efff34",
		16#082c# => X"e08c7805",
		16#082d# => X"e0632004",
		16#082e# => X"adef0030",
		16#082f# => X"e08d7805",
		16#0830# => X"e0632004",
		16#0831# => X"e08e7805",
		16#0832# => X"e0632004",
		16#0833# => X"d4401f04",
		16#0834# => X"18e00000",
		16#0835# => X"a8e71708",
		16#0836# => X"a880dead",
		16#0837# => X"dc402708",
		16#0838# => X"a8a0beef",
		16#0839# => X"dc072802",
		16#083a# => X"84c01708",
		16#083b# => X"1860dead",
		16#083c# => X"a863beef",
		16#083d# => X"e0633005",
		16#083e# => X"a9000012",
		16#083f# => X"d8404708",
		16#0840# => X"a9200034",
		16#0841# => X"d8074801",
		16#0842# => X"a9400056",
		16#0843# => X"d8075002",
		16#0844# => X"a9600078",
		16#0845# => X"d8075803",
		16#0846# => X"85870000",
		16#0847# => X"19a01234",
		16#0848# => X"a9ad5678",
		16#0849# => X"e1ad6005",
		16#084a# => X"e0636804",
		16#084b# => X"d4401f08",
		16#084c# => X"a800ffff",
		16#084d# => X"a8601234",
		16#084e# => X"9c832326",
		16#084f# => X"a0a3fcda",
		16#0850# => X"a0a5ffff",
		16#0851# => X"a4c32326",
		16#0852# => X"a8e32326",
		16#0853# => X"b1030005",
		16#0854# => X"b123fff5",
		16#0855# => X"e0243000",
		16#0856# => X"e0214000",
		16#0857# => X"9c219000",
		16#0858# => X"a021dd7d",
		16#0859# => X"e0453800",
		16#085a# => X"e0424800",
		16#085b# => X"a0427000",
		16#085c# => X"a04215f8",
		16#085d# => X"e0211004",
		16#085e# => X"d4400f0c",
		16#085f# => X"a9402326",
		16#0860# => X"a9600326",
		16#0861# => X"a9800005",
		16#0862# => X"ada0fff5",
		16#0863# => X"e1c35000",
		16#0864# => X"e1ce0001",
		16#0865# => X"e02e2005",
		16#0866# => X"e1c35802",
		16#0867# => X"e1ce0001",
		16#0868# => X"e04e2805",
		16#0869# => X"e0211004",
		16#086a# => X"e1c05002",
		16#086b# => X"a1ce2325",
		16#086c# => X"e0217004",
		16#086d# => X"e1c35003",
		16#086e# => X"e04e3005",
		16#086f# => X"e0211004",
		16#0870# => X"e1c35004",
		16#0871# => X"e04e3805",
		16#0872# => X"e0211004",
		16#0873# => X"e1c3630b",
		16#0874# => X"e04e4005",
		16#0875# => X"e0211004",
		16#0876# => X"e1c36b06",
		16#0877# => X"e04e4805",
		16#0878# => X"e0211004",
		16#0879# => X"d4400f10",
		16#087a# => X"ac60ffff",
		16#087b# => X"9c230001",
		16#087c# => X"a483ffff",
		16#087d# => X"a8a4ffff",
		16#087e# => X"9cc58000",
		16#087f# => X"ac467fff",
		16#0880# => X"e0211004",
		16#0881# => X"b0e3ffff",
		16#0882# => X"ac470001",
		16#0883# => X"e0211004",
		16#0884# => X"d4400f14",
		16#0885# => X"a8200001",
		16#0886# => X"a840000a",
		16#0887# => X"a8600015",
		16#0888# => X"18804040",
		16#0889# => X"a8841010",
		16#088a# => X"e0a40808",
		16#088b# => X"e0c11008",
		16#088c# => X"e0e11808",
		16#088d# => X"e1040848",
		16#088e# => X"e1251048",
		16#088f# => X"e1451848",
		16#0890# => X"e1640888",
		16#0891# => X"e1851088",
		16#0892# => X"e1a51888",
		16#0893# => X"e0253005",
		16#0894# => X"e0474005",
		16#0895# => X"e0695005",
		16#0896# => X"e08b6005",
		16#0897# => X"e0216805",
		16#0898# => X"e0421805",
		16#0899# => X"e0212005",
		16#089a# => X"e0211005",
		16#089b# => X"1840809f",
		16#089c# => X"a842dc20",
		16#089d# => X"e0211005",
		16#089e# => X"d4400f18",
		16#089f# => X"a8200001",
		16#08a0# => X"ac60fffb",
		16#08a1# => X"a8400001",
		16#08a2# => X"e4011800",
		16#08a3# => X"e082000e",
		16#08a4# => X"e0a02004",
		16#08a5# => X"e4030800",
		16#08a6# => X"e082000e",
		16#08a7# => X"e0a52004",
		16#08a8# => X"e4021000",
		16#08a9# => X"e080100e",
		16#08aa# => X"e0a52004",
		16#08ab# => X"a8400002",
		16#08ac# => X"e4211800",
		16#08ad# => X"e080100e",
		16#08ae# => X"e0a52004",
		16#08af# => X"e4230800",
		16#08b0# => X"e080100e",
		16#08b1# => X"e0a52004",
		16#08b2# => X"e4221000",
		16#08b3# => X"e082000e",
		16#08b4# => X"e0a52004",
		16#08b5# => X"a8400004",
		16#08b6# => X"e4411800",
		16#08b7# => X"e082000e",
		16#08b8# => X"e0a52004",
		16#08b9# => X"e4430800",
		16#08ba# => X"e080100e",
		16#08bb# => X"e0a52004",
		16#08bc# => X"e4421000",
		16#08bd# => X"e082000e",
		16#08be# => X"e0a52004",
		16#08bf# => X"a8400008",
		16#08c0# => X"e4611800",
		16#08c1# => X"e082000e",
		16#08c2# => X"e0a52004",
		16#08c3# => X"e4630800",
		16#08c4# => X"e080100e",
		16#08c5# => X"e0a52004",
		16#08c6# => X"e4621000",
		16#08c7# => X"e080100e",
		16#08c8# => X"e0a52004",
		16#08c9# => X"a8400010",
		16#08ca# => X"e4811800",
		16#08cb# => X"e080100e",
		16#08cc# => X"e0a52004",
		16#08cd# => X"e4830800",
		16#08ce# => X"e082000e",
		16#08cf# => X"e0a52004",
		16#08d0# => X"e4821000",
		16#08d1# => X"e082000e",
		16#08d2# => X"e0a52004",
		16#08d3# => X"a8400020",
		16#08d4# => X"e4a11800",
		16#08d5# => X"e080100e",
		16#08d6# => X"e0a52004",
		16#08d7# => X"e4a30800",
		16#08d8# => X"e082000e",
		16#08d9# => X"e0a52004",
		16#08da# => X"e4a21000",
		16#08db# => X"e080100e",
		16#08dc# => X"e0a52004",
		16#08dd# => X"a8400040",
		16#08de# => X"e5411800",
		16#08df# => X"e080100e",
		16#08e0# => X"e0a52004",
		16#08e1# => X"e5430800",
		16#08e2# => X"e082000e",
		16#08e3# => X"e0a52004",
		16#08e4# => X"e5400800",
		16#08e5# => X"e082000e",
		16#08e6# => X"e0a52004",
		16#08e7# => X"e5410000",
		16#08e8# => X"e080100e",
		16#08e9# => X"e0a52004",
		16#08ea# => X"e5421000",
		16#08eb# => X"e082000e",
		16#08ec# => X"e0a52004",
		16#08ed# => X"a8400080",
		16#08ee# => X"e5611800",
		16#08ef# => X"e080100e",
		16#08f0# => X"e0a52004",
		16#08f1# => X"e5630800",
		16#08f2# => X"e082000e",
		16#08f3# => X"e0a52004",
		16#08f4# => X"e5600800",
		16#08f5# => X"e082000e",
		16#08f6# => X"e0a52004",
		16#08f7# => X"e5610000",
		16#08f8# => X"e080100e",
		16#08f9# => X"e0a52004",
		16#08fa# => X"e5621000",
		16#08fb# => X"e080100e",
		16#08fc# => X"e0a52004",
		16#08fd# => X"a8400100",
		16#08fe# => X"e5811800",
		16#08ff# => X"e082000e",
		16#0900# => X"e0a52004",
		16#0901# => X"e5830800",
		16#0902# => X"e080100e",
		16#0903# => X"e0a52004",
		16#0904# => X"e5800800",
		16#0905# => X"e080100e",
		16#0906# => X"e0a52004",
		16#0907# => X"e5810000",
		16#0908# => X"e082000e",
		16#0909# => X"e0a52004",
		16#090a# => X"e5821000",
		16#090b# => X"e082000e",
		16#090c# => X"e0a52004",
		16#090d# => X"a8400200",
		16#090e# => X"e5a11800",
		16#090f# => X"e082000e",
		16#0910# => X"e0a52004",
		16#0911# => X"e5a30800",
		16#0912# => X"e080100e",
		16#0913# => X"e0a52004",
		16#0914# => X"e5a00800",
		16#0915# => X"e080100e",
		16#0916# => X"e0a52004",
		16#0917# => X"e5a10000",
		16#0918# => X"e082000e",
		16#0919# => X"e0a52004",
		16#091a# => X"e5a21000",
		16#091b# => X"e080100e",
		16#091c# => X"e0a52004",
		16#091d# => X"d4402f1c",
		16#091e# => X"a8200011",
		16#091f# => X"ac60fff7",
		16#0920# => X"a8400001",
		16#0921# => X"bc01fff7",
		16#0922# => X"e082000e",
		16#0923# => X"e0a02004",
		16#0924# => X"bc030011",
		16#0925# => X"e082000e",
		16#0926# => X"e0a52004",
		16#0927# => X"bc010011",
		16#0928# => X"e080100e",
		16#0929# => X"e0a52004",
		16#092a# => X"a8400002",
		16#092b# => X"bc21fff7",
		16#092c# => X"e080100e",
		16#092d# => X"e0a52004",
		16#092e# => X"bc230011",
		16#092f# => X"e080100e",
		16#0930# => X"e0a52004",
		16#0931# => X"bc210011",
		16#0932# => X"e082000e",
		16#0933# => X"e0a52004",
		16#0934# => X"a8400004",
		16#0935# => X"bc41fff7",
		16#0936# => X"e082000e",
		16#0937# => X"e0a52004",
		16#0938# => X"bc430011",
		16#0939# => X"e080100e",
		16#093a# => X"e0a52004",
		16#093b# => X"bc410011",
		16#093c# => X"e082000e",
		16#093d# => X"e0a52004",
		16#093e# => X"a8400008",
		16#093f# => X"bc61fff7",
		16#0940# => X"e082000e",
		16#0941# => X"e0a52004",
		16#0942# => X"bc630011",
		16#0943# => X"e080100e",
		16#0944# => X"e0a52004",
		16#0945# => X"bc610011",
		16#0946# => X"e080100e",
		16#0947# => X"e0a52004",
		16#0948# => X"a8400010",
		16#0949# => X"bc81fff7",
		16#094a# => X"e080100e",
		16#094b# => X"e0a52004",
		16#094c# => X"bc830011",
		16#094d# => X"e082000e",
		16#094e# => X"e0a52004",
		16#094f# => X"bc810011",
		16#0950# => X"e082000e",
		16#0951# => X"e0a52004",
		16#0952# => X"a8400020",
		16#0953# => X"bca1fff7",
		16#0954# => X"e080100e",
		16#0955# => X"e0a52004",
		16#0956# => X"bca30011",
		16#0957# => X"e082000e",
		16#0958# => X"e0a52004",
		16#0959# => X"bca10011",
		16#095a# => X"e080100e",
		16#095b# => X"e0a52004",
		16#095c# => X"a8400040",
		16#095d# => X"bd41fff7",
		16#095e# => X"e080100e",
		16#095f# => X"e0a52004",
		16#0960# => X"bd430011",
		16#0961# => X"e082000e",
		16#0962# => X"e0a52004",
		16#0963# => X"bd400011",
		16#0964# => X"e082000e",
		16#0965# => X"e0a52004",
		16#0966# => X"bd410000",
		16#0967# => X"e080100e",
		16#0968# => X"e0a52004",
		16#0969# => X"bd410011",
		16#096a# => X"e082000e",
		16#096b# => X"e0a52004",
		16#096c# => X"a8400080",
		16#096d# => X"bd61fff7",
		16#096e# => X"e080100e",
		16#096f# => X"e0a52004",
		16#0970# => X"bd630011",
		16#0971# => X"e082000e",
		16#0972# => X"e0a52004",
		16#0973# => X"bd600011",
		16#0974# => X"e082000e",
		16#0975# => X"e0a52004",
		16#0976# => X"bd610000",
		16#0977# => X"e080100e",
		16#0978# => X"e0a52004",
		16#0979# => X"bd610011",
		16#097a# => X"e080100e",
		16#097b# => X"e0a52004",
		16#097c# => X"a8400100",
		16#097d# => X"bd81fff7",
		16#097e# => X"e082000e",
		16#097f# => X"e0a52004",
		16#0980# => X"bd830011",
		16#0981# => X"e080100e",
		16#0982# => X"e0a52004",
		16#0983# => X"bd800011",
		16#0984# => X"e080100e",
		16#0985# => X"e0a52004",
		16#0986# => X"bd810000",
		16#0987# => X"e082000e",
		16#0988# => X"e0a52004",
		16#0989# => X"bd810011",
		16#098a# => X"e082000e",
		16#098b# => X"e0a52004",
		16#098c# => X"a8400200",
		16#098d# => X"bda1fff7",
		16#098e# => X"e082000e",
		16#098f# => X"e0a52004",
		16#0990# => X"bda30011",
		16#0991# => X"e080100e",
		16#0992# => X"e0a52004",
		16#0993# => X"bda00011",
		16#0994# => X"e080100e",
		16#0995# => X"e0a52004",
		16#0996# => X"bda10000",
		16#0997# => X"e082000e",
		16#0998# => X"e0a52004",
		16#0999# => X"bda10011",
		16#099a# => X"e080100e",
		16#099b# => X"e0a52004",
		16#099c# => X"d4402f20",
		16#099d# => X"15000000",
		16#099e# => X"a8200001",
		16#099f# => X"00000006",
		16#09a0# => X"ac210001",
		16#09a1# => X"a8210001",
		16#09a2# => X"e0400004",
		16#09a3# => X"00000005",
		16#09a4# => X"15000000",
		16#09a5# => X"a8400001",
		16#09a6# => X"03fffffc",
		16#09a7# => X"15000000",
		16#09a8# => X"e0211004",
		16#09a9# => X"a8400002",
		16#09aa# => X"a86026b8",
		16#09ab# => X"44001800",
		16#09ac# => X"ac420002",
		16#09ad# => X"a8420002",
		16#09ae# => X"e0211004",
		16#09af# => X"a8400004",
		16#09b0# => X"04000003",
		16#09b1# => X"ac420004",
		16#09b2# => X"a8420004",
		16#09b3# => X"a86026c8",
		16#09b4# => X"a8800004",
		16#09b5# => X"e4034800",
		16#09b6# => X"e042200e",
		16#09b7# => X"e0211004",
		16#09b8# => X"a8400008",
		16#09b9# => X"a86026f4",
		16#09ba# => X"48001800",
		16#09bb# => X"ac420008",
		16#09bc# => X"a8420008",
		16#09bd# => X"a86026f0",
		16#09be# => X"a8800008",
		16#09bf# => X"e4034800",
		16#09c0# => X"e042200e",
		16#09c1# => X"e0211004",
		16#09c2# => X"a84000f0",
		16#09c3# => X"e4000000",
		16#09c4# => X"10000003",
		16#09c5# => X"ac420010",
		16#09c6# => X"a8420010",
		16#09c7# => X"0c000003",
		16#09c8# => X"15000000",
		16#09c9# => X"ac420080",
		16#09ca# => X"e4200000",
		16#09cb# => X"0c000003",
		16#09cc# => X"ac420040",
		16#09cd# => X"a8420040",
		16#09ce# => X"10000003",
		16#09cf# => X"15000000",
		16#09d0# => X"ac420020",
		16#09d1# => X"e0211004",
		16#09d2# => X"d4400f24",
		16#09d3# => X"15000001",
		16#09d4# => X"00000000",
		others => X"00000000"
	);

end package;