library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.types.all;

package prog_mem is

	constant PROG_SIZE : integer := 8268;

	constant PROG_DATA : mem_type(0 to PROG_SIZE/4-1) := (
		16#0000# => X"97100000",
		16#0001# => X"93800000",
		16#0002# => X"73905030",
		16#0003# => X"f32040f1",
		16#0004# => X"63860000",
		16#0005# => X"f090f090",
		16#0006# => X"0b000000",
		16#0007# => X"97200000",
		16#0008# => X"938040fe",
		16#0009# => X"37c1feca",
		16#000a# => X"1301e1ab",
		16#000b# => X"23a02000",
		16#000c# => X"0bb00000",
		16#000d# => X"83a10000",
		16#000e# => X"631c3178",
		16#000f# => X"97270000",
		16#0010# => X"938707ff",
		16#0011# => X"37c7adde",
		16#0012# => X"1307f7ee",
		16#0013# => X"83a60700",
		16#0014# => X"6390e678",
		16#0015# => X"1301e0fb",
		16#0016# => X"83810000",
		16#0017# => X"1302a0fb",
		16#0018# => X"83821000",
		16#0019# => X"1303e0ff",
		16#001a# => X"83832000",
		16#001b# => X"1304a0fc",
		16#001c# => X"83843000",
		16#001d# => X"631e3174",
		16#001e# => X"631c5274",
		16#001f# => X"631a7374",
		16#0020# => X"63189474",
		16#0021# => X"37c1ffff",
		16#0022# => X"1301e1ab",
		16#0023# => X"83910000",
		16#0024# => X"37d2ffff",
		16#0025# => X"1302e2af",
		16#0026# => X"83922000",
		16#0027# => X"631a3172",
		16#0028# => X"63185272",
		16#0029# => X"37c10000",
		16#002a# => X"1301e1ab",
		16#002b# => X"83d10000",
		16#002c# => X"37d20000",
		16#002d# => X"1302e2af",
		16#002e# => X"83d22000",
		16#002f# => X"631a3170",
		16#0030# => X"63185270",
		16#0031# => X"1301e00b",
		16#0032# => X"83c10000",
		16#0033# => X"1302a00b",
		16#0034# => X"83c21000",
		16#0035# => X"1303e00f",
		16#0036# => X"83c32000",
		16#0037# => X"1304a00c",
		16#0038# => X"83c43000",
		16#0039# => X"6316316e",
		16#003a# => X"6314526e",
		16#003b# => X"6312736e",
		16#003c# => X"6310946e",
		16#003d# => X"97200000",
		16#003e# => X"938000f5",
		16#003f# => X"37d10000",
		16#0040# => X"1301e1af",
		16#0041# => X"b7c10000",
		16#0042# => X"9381e1ab",
		16#0043# => X"b7c2feca",
		16#0044# => X"9382e2ab",
		16#0045# => X"23912000",
		16#0046# => X"0bb00000",
		16#0047# => X"23903000",
		16#0048# => X"0bb00000",
		16#0049# => X"03d22000",
		16#004a# => X"6314416a",
		16#004b# => X"03d20000",
		16#004c# => X"6390416a",
		16#004d# => X"03a20000",
		16#004e# => X"639c4268",
		16#004f# => X"1301500a",
		16#0050# => X"b7a2a3a2",
		16#0051# => X"9382524a",
		16#0052# => X"23802000",
		16#0053# => X"03c20000",
		16#0054# => X"63104168",
		16#0055# => X"1301f1ff",
		16#0056# => X"a3802000",
		16#0057# => X"03c21000",
		16#0058# => X"63184166",
		16#0059# => X"1301f1ff",
		16#005a# => X"23812000",
		16#005b# => X"03c22000",
		16#005c# => X"63104166",
		16#005d# => X"1301f1ff",
		16#005e# => X"a3812000",
		16#005f# => X"03c23000",
		16#0060# => X"63184164",
		16#0061# => X"83a10000",
		16#0062# => X"63945164",
		16#0063# => X"97200000",
		16#0064# => X"938080e7",
		16#0065# => X"17210000",
		16#0066# => X"130141e7",
		16#0067# => X"23a00000",
		16#0068# => X"23200100",
		16#0069# => X"13000000",
		16#006a# => X"972f0000",
		16#006b# => X"938f4fe6",
		16#006c# => X"370f0090",
		16#006d# => X"93004006",
		16#006e# => X"23201f00",
		16#006f# => X"93003012",
		16#0070# => X"9380d0dd",
		16#0071# => X"93800010",
		16#0072# => X"23801f00",
		16#0073# => X"1360f07f",
		16#0074# => X"93e03012",
		16#0075# => X"93e01032",
		16#0076# => X"1381d0cd",
		16#0077# => X"a3802f00",
		16#0078# => X"93f0007f",
		16#0079# => X"93f0f07f",
		16#007a# => X"138100ce",
		16#007b# => X"23812f00",
		16#007c# => X"93c05075",
		16#007d# => X"93c05047",
		16#007e# => X"a3811f00",
		16#007f# => X"83a00f00",
		16#0080# => X"6318105c",
		16#0081# => X"13000000",
		16#0082# => X"972f0000",
		16#0083# => X"938f8fe0",
		16#0084# => X"b7a0a5a5",
		16#0085# => X"9380505a",
		16#0086# => X"37c1feca",
		16#0087# => X"1301e1ab",
		16#0088# => X"b701feca",
		16#0089# => X"37c20000",
		16#008a# => X"1302e2ab",
		16#008b# => X"b7c20000",
		16#008c# => X"9382f2ee",
		16#008d# => X"b7a25b6f",
		16#008e# => X"9382525a",
		16#008f# => X"13653012",
		16#0090# => X"93656024",
		16#0091# => X"3306b540",
		16#0092# => X"3306a600",
		16#0093# => X"2380cf00",
		16#0094# => X"33e54100",
		16#0095# => X"b3052540",
		16#0096# => X"a380bf00",
		16#0097# => X"b3753500",
		16#0098# => X"b3853540",
		16#0099# => X"2381bf00",
		16#009a# => X"b3454500",
		16#009b# => X"b3c51500",
		16#009c# => X"b3c55500",
		16#009d# => X"a381bf00",
		16#009e# => X"83a00f00",
		16#009f# => X"631a1054",
		16#00a0# => X"13000000",
		16#00a1# => X"972f0000",
		16#00a2# => X"938f0fd9",
		16#00a3# => X"93001000",
		16#00a4# => X"1301a000",
		16#00a5# => X"93015001",
		16#00a6# => X"37124040",
		16#00a7# => X"13020201",
		16#00a8# => X"b3120200",
		16#00a9# => X"33530200",
		16#00aa# => X"b3530240",
		16#00ab# => X"33c46200",
		16#00ac# => X"b3447200",
		16#00ad# => X"33659400",
		16#00ae# => X"2380af00",
		16#00af# => X"631a0550",
		16#00b0# => X"b3121200",
		16#00b1# => X"33932000",
		16#00b2# => X"b3933000",
		16#00b3# => X"33541200",
		16#00b4# => X"b3d42200",
		16#00b5# => X"33d53200",
		16#00b6# => X"b3551240",
		16#00b7# => X"33d62240",
		16#00b8# => X"b3d63240",
		16#00b9# => X"b3c06200",
		16#00ba# => X"33c18300",
		16#00bb# => X"b3c1a400",
		16#00bc# => X"33c2c500",
		16#00bd# => X"b3c0d000",
		16#00be# => X"33413100",
		16#00bf# => X"b3c04000",
		16#00c0# => X"b3c02000",
		16#00c1# => X"37e19f80",
		16#00c2# => X"130101c2",
		16#00c3# => X"b3c02000",
		16#00c4# => X"a3801f00",
		16#00c5# => X"93001000",
		16#00c6# => X"1301a000",
		16#00c7# => X"93015001",
		16#00c8# => X"37124040",
		16#00c9# => X"13020201",
		16#00ca# => X"93121200",
		16#00cb# => X"1393a000",
		16#00cc# => X"93935001",
		16#00cd# => X"13541200",
		16#00ce# => X"93d4a200",
		16#00cf# => X"13d55201",
		16#00d0# => X"93551240",
		16#00d1# => X"13d6a240",
		16#00d2# => X"93d65241",
		16#00d3# => X"b3c06200",
		16#00d4# => X"33c18300",
		16#00d5# => X"b3c1a400",
		16#00d6# => X"33c2c500",
		16#00d7# => X"b3c0d000",
		16#00d8# => X"33413100",
		16#00d9# => X"b3c04000",
		16#00da# => X"b3c02000",
		16#00db# => X"37e19f80",
		16#00dc# => X"130101c2",
		16#00dd# => X"b3c02000",
		16#00de# => X"23911f00",
		16#00df# => X"83a00f00",
		16#00e0# => X"63181044",
		16#00e1# => X"13000000",
		16#00e2# => X"972f0000",
		16#00e3# => X"938f0fc9",
		16#00e4# => X"93002003",
		16#00e5# => X"1301e0fc",
		16#00e6# => X"9303b007",
		16#00e7# => X"130450f8",
		16#00e8# => X"93041000",
		16#00e9# => X"1305f0ff",
		16#00ea# => X"93a1b007",
		16#00eb# => X"13a250f8",
		16#00ec# => X"9322b107",
		16#00ed# => X"132351f8",
		16#00ee# => X"b3c15100",
		16#00ef# => X"33426200",
		16#00f0# => X"b3e54100",
		16#00f1# => X"2380bf00",
		16#00f2# => X"93b150f8",
		16#00f3# => X"13b21000",
		16#00f4# => X"9332f1ff",
		16#00f5# => X"1333b107",
		16#00f6# => X"b3c15100",
		16#00f7# => X"33426200",
		16#00f8# => X"b3e54100",
		16#00f9# => X"a380bf00",
		16#00fa# => X"b3a17000",
		16#00fb# => X"33a28000",
		16#00fc# => X"b3227100",
		16#00fd# => X"33238100",
		16#00fe# => X"b3c15100",
		16#00ff# => X"33426200",
		16#0100# => X"b3e54100",
		16#0101# => X"2381bf00",
		16#0102# => X"b3b18000",
		16#0103# => X"33b29000",
		16#0104# => X"b332a100",
		16#0105# => X"33337100",
		16#0106# => X"b3c15100",
		16#0107# => X"33426200",
		16#0108# => X"b3e54100",
		16#0109# => X"a381bf00",
		16#010a# => X"83a00f00",
		16#010b# => X"6312103a",
		16#010c# => X"13000000",
		16#010d# => X"972f0000",
		16#010e# => X"938f8fbe",
		16#010f# => X"13000000",
		16#0110# => X"13000000",
		16#0111# => X"b3600000",
		16#0112# => X"6f004001",
		16#0113# => X"93e01000",
		16#0114# => X"13411100",
		16#0115# => X"6f000001",
		16#0116# => X"13000000",
		16#0117# => X"13611000",
		16#0118# => X"6ff01fff",
		16#0119# => X"b3e02000",
		16#011a# => X"13610000",
		16#011b# => X"97010000",
		16#011c# => X"93810101",
		16#011d# => X"67800100",
		16#011e# => X"13612100",
		16#011f# => X"b3e02000",
		16#0120# => X"33610000",
		16#0121# => X"ef048000",
		16#0122# => X"13614100",
		16#0123# => X"97010000",
		16#0124# => X"9381c1ff",
		16#0125# => X"b3c19100",
		16#0126# => X"b3e02000",
		16#0127# => X"b3e03000",
		16#0128# => X"33610000",
		16#0129# => X"97010000",
		16#012a# => X"93810101",
		16#012b# => X"e7840100",
		16#012c# => X"13618100",
		16#012d# => X"97010000",
		16#012e# => X"9381c1ff",
		16#012f# => X"b3c19100",
		16#0130# => X"b3e02000",
		16#0131# => X"b3e03000",
		16#0132# => X"23901f00",
		16#0133# => X"13010000",
		16#0134# => X"93012003",
		16#0135# => X"1302e0fc",
		16#0136# => X"93024006",
		16#0137# => X"1303c0f9",
		16#0138# => X"93031000",
		16#0139# => X"1304f0ff",
		16#013a# => X"13056009",
		16#013b# => X"6302712e",
		16#013c# => X"33417100",
		16#013d# => X"63167100",
		16#013e# => X"e30c71fe",
		16#013f# => X"13612100",
		16#0140# => X"33053540",
		16#0141# => X"e34ea4fe",
		16#0142# => X"33057500",
		16#0143# => X"e35ea4fe",
		16#0144# => X"3361a100",
		16#0145# => X"33057500",
		16#0146# => X"e36e35fe",
		16#0147# => X"33057540",
		16#0148# => X"e37e85fe",
		16#0149# => X"13051500",
		16#014a# => X"33453500",
		16#014b# => X"3361a100",
		16#014c# => X"23912f00",
		16#014d# => X"03a10f00",
		16#014e# => X"631c2028",
		16#014f# => X"972f0000",
		16#0150# => X"938f4fae",
		16#0151# => X"97100000",
		16#0152# => X"9380c0ab",
		16#0153# => X"73905030",
		16#0154# => X"93000000",
		16#0155# => X"13013000",
		16#0156# => X"93801000",
		16#0157# => X"f090f090",
		16#0158# => X"93802000",
		16#0159# => X"b3c02000",
		16#015a# => X"23801f00",
		16#015b# => X"93008008",
		16#015c# => X"1301f0ff",
		16#015d# => X"93010000",
		16#015e# => X"731510f1",
		16#015f# => X"73900030",
		16#0160# => X"f3250030",
		16#0161# => X"73100130",
		16#0162# => X"73260030",
		16#0163# => X"33cec500",
		16#0164# => X"b34e3500",
		16#0165# => X"336fc001",
		16#0166# => X"336fdf01",
		16#0167# => X"733510f1",
		16#0168# => X"733511f1",
		16#0169# => X"73b00030",
		16#016a# => X"f3250030",
		16#016b# => X"73300130",
		16#016c# => X"73260030",
		16#016d# => X"33cec500",
		16#016e# => X"b34e3500",
		16#016f# => X"336fcf01",
		16#0170# => X"336fdf01",
		16#0171# => X"a380ef01",
		16#0172# => X"735510f1",
		16#0173# => X"73500430",
		16#0174# => X"f3250030",
		16#0175# => X"73d00f30",
		16#0176# => X"73260030",
		16#0177# => X"33cec500",
		16#0178# => X"b34e3500",
		16#0179# => X"336fcf01",
		16#017a# => X"336fdf01",
		16#017b# => X"737510f1",
		16#017c# => X"73f51ff1",
		16#017d# => X"73700430",
		16#017e# => X"f3250030",
		16#017f# => X"73f00f30",
		16#0180# => X"73260030",
		16#0181# => X"33cec500",
		16#0182# => X"b34e3500",
		16#0183# => X"336fcf01",
		16#0184# => X"336fdf01",
		16#0185# => X"2381ef01",
		16#0186# => X"732510f1",
		16#0187# => X"732511f1",
		16#0188# => X"73a00030",
		16#0189# => X"f3250030",
		16#018a# => X"73200130",
		16#018b# => X"73260030",
		16#018c# => X"33cec500",
		16#018d# => X"b34e3500",
		16#018e# => X"336fcf01",
		16#018f# => X"336fdf01",
		16#0190# => X"736510f1",
		16#0191# => X"73e51ff1",
		16#0192# => X"73600430",
		16#0193# => X"f3250030",
		16#0194# => X"73e00f30",
		16#0195# => X"73260030",
		16#0196# => X"33cec500",
		16#0197# => X"b34e3500",
		16#0198# => X"336fcf01",
		16#0199# => X"336fdf01",
		16#019a# => X"a381ef01",
		16#019b# => X"93007000",
		16#019c# => X"17210000",
		16#019d# => X"1301019c",
		16#019e# => X"03210100",
		16#019f# => X"639a2014",
		16#01a0# => X"83a10f00",
		16#01a1# => X"63960114",
		16#01a2# => X"972f0000",
		16#01a3# => X"938fcf99",
		16#01a4# => X"172f0000",
		16#01a5# => X"130f4f9a",
		16#01a6# => X"83a01f00",
		16#01a7# => X"83a02f00",
		16#01a8# => X"83a03f00",
		16#01a9# => X"83901f00",
		16#01aa# => X"83903f00",
		16#01ab# => X"03210f00",
		16#01ac# => X"93405100",
		16#01ad# => X"23801f00",
		16#01ae# => X"172f0000",
		16#01af# => X"130f0f98",
		16#01b0# => X"b7c0feca",
		16#01b1# => X"9380e0ab",
		16#01b2# => X"a3a01f00",
		16#01b3# => X"23a11f00",
		16#01b4# => X"a3a11f00",
		16#01b5# => X"a3901f00",
		16#01b6# => X"a3911f00",
		16#01b7# => X"03210f00",
		16#01b8# => X"93405100",
		16#01b9# => X"a3801f00",
		16#01ba# => X"172f0000",
		16#01bb# => X"130f4f95",
		16#01bc# => X"97000000",
		16#01bd# => X"9380000e",
		16#01be# => X"6f002000",
		16#01bf# => X"67802000",
		16#01c0# => X"6780f01f",
		16#01c1# => X"63010000",
		16#01c2# => X"e31f1000",
		16#01c3# => X"e34f1000",
		16#01c4# => X"63041000",
		16#01c5# => X"03210f00",
		16#01c6# => X"93406100",
		16#01c7# => X"23811f00",
		16#01c8# => X"a3811f00",
		16#01c9# => X"83a10f00",
		16#01ca# => X"972f0000",
		16#01cb# => X"938f0f90",
		16#01cc# => X"73211030",
		16#01cd# => X"b7110000",
		16#01ce# => X"b3713100",
		16#01cf# => X"638a0106",
		16#01d0# => X"93002000",
		16#01d1# => X"13015000",
		16#01d2# => X"9301a000",
		16#01d3# => X"37a29999",
		16#01d4# => X"13029299",
		16#01d5# => X"9302d0ff",
		16#01d6# => X"1303f0ff",
		16#01d7# => X"b3832002",
		16#01d8# => X"b3833302",
		16#01d9# => X"b3831302",
		16#01da# => X"93c3830c",
		16#01db# => X"63127006",
		16#01dc# => X"b3836002",
		16#01dd# => X"b3833302",
		16#01de# => X"b3835302",
		16#01df# => X"93c3c303",
		16#01e0# => X"63187004",
		16#01e1# => X"b3834002",
		16#01e2# => X"b3934002",
		16#01e3# => X"73001000",
		16#01e4# => X"93001000",
		16#01e5# => X"b3231302",
		16#01e6# => X"b3c32102",
		16#01e7# => X"b3433102",
		16#01e8# => X"b3e32102",
		16#01e9# => X"b3633102",
		16#01ea# => X"23800f00",
		16#01eb# => X"6f00c000",
		16#01ec# => X"9300a00a",
		16#01ed# => X"23801f00",
		16#01ee# => X"9300b00b",
		16#01ef# => X"a3801f00",
		16#01f0# => X"9300c00c",
		16#01f1# => X"23811f00",
		16#01f2# => X"9300d00d",
		16#01f3# => X"a3811f00",
		16#01f4# => X"97200000",
		16#01f5# => X"93800083",
		16#01f6# => X"0bb00000",
		16#01f7# => X"0b000000",
		16#01f8# => X"00000000",
		16#01f9# => X"00000000",
		16#01fa# => X"00000000",
		16#01fb# => X"00000000",
		16#01fc# => X"00000000",
		16#01fd# => X"00000000",
		16#01fe# => X"00000000",
		16#01ff# => X"00000000",
		16#0200# => X"00000000",
		16#0201# => X"00000000",
		16#0202# => X"00000000",
		16#0203# => X"00000000",
		16#0204# => X"00000000",
		16#0205# => X"00000000",
		16#0206# => X"00000000",
		16#0207# => X"00000000",
		16#0208# => X"00000000",
		16#0209# => X"00000000",
		16#020a# => X"00000000",
		16#020b# => X"00000000",
		16#020c# => X"00000000",
		16#020d# => X"00000000",
		16#020e# => X"00000000",
		16#020f# => X"00000000",
		16#0210# => X"00000000",
		16#0211# => X"00000000",
		16#0212# => X"00000000",
		16#0213# => X"00000000",
		16#0214# => X"00000000",
		16#0215# => X"00000000",
		16#0216# => X"00000000",
		16#0217# => X"00000000",
		16#0218# => X"00000000",
		16#0219# => X"00000000",
		16#021a# => X"00000000",
		16#021b# => X"00000000",
		16#021c# => X"00000000",
		16#021d# => X"00000000",
		16#021e# => X"00000000",
		16#021f# => X"00000000",
		16#0220# => X"00000000",
		16#0221# => X"00000000",
		16#0222# => X"00000000",
		16#0223# => X"00000000",
		16#0224# => X"00000000",
		16#0225# => X"00000000",
		16#0226# => X"00000000",
		16#0227# => X"00000000",
		16#0228# => X"00000000",
		16#0229# => X"00000000",
		16#022a# => X"00000000",
		16#022b# => X"00000000",
		16#022c# => X"00000000",
		16#022d# => X"00000000",
		16#022e# => X"00000000",
		16#022f# => X"00000000",
		16#0230# => X"00000000",
		16#0231# => X"00000000",
		16#0232# => X"00000000",
		16#0233# => X"00000000",
		16#0234# => X"00000000",
		16#0235# => X"00000000",
		16#0236# => X"00000000",
		16#0237# => X"00000000",
		16#0238# => X"00000000",
		16#0239# => X"00000000",
		16#023a# => X"00000000",
		16#023b# => X"00000000",
		16#023c# => X"00000000",
		16#023d# => X"00000000",
		16#023e# => X"00000000",
		16#023f# => X"00000000",
		16#0240# => X"00000000",
		16#0241# => X"00000000",
		16#0242# => X"00000000",
		16#0243# => X"00000000",
		16#0244# => X"00000000",
		16#0245# => X"00000000",
		16#0246# => X"00000000",
		16#0247# => X"00000000",
		16#0248# => X"00000000",
		16#0249# => X"00000000",
		16#024a# => X"00000000",
		16#024b# => X"00000000",
		16#024c# => X"00000000",
		16#024d# => X"00000000",
		16#024e# => X"00000000",
		16#024f# => X"00000000",
		16#0250# => X"00000000",
		16#0251# => X"00000000",
		16#0252# => X"00000000",
		16#0253# => X"00000000",
		16#0254# => X"00000000",
		16#0255# => X"00000000",
		16#0256# => X"00000000",
		16#0257# => X"00000000",
		16#0258# => X"00000000",
		16#0259# => X"00000000",
		16#025a# => X"00000000",
		16#025b# => X"00000000",
		16#025c# => X"00000000",
		16#025d# => X"00000000",
		16#025e# => X"00000000",
		16#025f# => X"00000000",
		16#0260# => X"00000000",
		16#0261# => X"00000000",
		16#0262# => X"00000000",
		16#0263# => X"00000000",
		16#0264# => X"00000000",
		16#0265# => X"00000000",
		16#0266# => X"00000000",
		16#0267# => X"00000000",
		16#0268# => X"00000000",
		16#0269# => X"00000000",
		16#026a# => X"00000000",
		16#026b# => X"00000000",
		16#026c# => X"00000000",
		16#026d# => X"00000000",
		16#026e# => X"00000000",
		16#026f# => X"00000000",
		16#0270# => X"00000000",
		16#0271# => X"00000000",
		16#0272# => X"00000000",
		16#0273# => X"00000000",
		16#0274# => X"00000000",
		16#0275# => X"00000000",
		16#0276# => X"00000000",
		16#0277# => X"00000000",
		16#0278# => X"00000000",
		16#0279# => X"00000000",
		16#027a# => X"00000000",
		16#027b# => X"00000000",
		16#027c# => X"00000000",
		16#027d# => X"00000000",
		16#027e# => X"00000000",
		16#027f# => X"00000000",
		16#0280# => X"00000000",
		16#0281# => X"00000000",
		16#0282# => X"00000000",
		16#0283# => X"00000000",
		16#0284# => X"00000000",
		16#0285# => X"00000000",
		16#0286# => X"00000000",
		16#0287# => X"00000000",
		16#0288# => X"00000000",
		16#0289# => X"00000000",
		16#028a# => X"00000000",
		16#028b# => X"00000000",
		16#028c# => X"00000000",
		16#028d# => X"00000000",
		16#028e# => X"00000000",
		16#028f# => X"00000000",
		16#0290# => X"00000000",
		16#0291# => X"00000000",
		16#0292# => X"00000000",
		16#0293# => X"00000000",
		16#0294# => X"00000000",
		16#0295# => X"00000000",
		16#0296# => X"00000000",
		16#0297# => X"00000000",
		16#0298# => X"00000000",
		16#0299# => X"00000000",
		16#029a# => X"00000000",
		16#029b# => X"00000000",
		16#029c# => X"00000000",
		16#029d# => X"00000000",
		16#029e# => X"00000000",
		16#029f# => X"00000000",
		16#02a0# => X"00000000",
		16#02a1# => X"00000000",
		16#02a2# => X"00000000",
		16#02a3# => X"00000000",
		16#02a4# => X"00000000",
		16#02a5# => X"00000000",
		16#02a6# => X"00000000",
		16#02a7# => X"00000000",
		16#02a8# => X"00000000",
		16#02a9# => X"00000000",
		16#02aa# => X"00000000",
		16#02ab# => X"00000000",
		16#02ac# => X"00000000",
		16#02ad# => X"00000000",
		16#02ae# => X"00000000",
		16#02af# => X"00000000",
		16#02b0# => X"00000000",
		16#02b1# => X"00000000",
		16#02b2# => X"00000000",
		16#02b3# => X"00000000",
		16#02b4# => X"00000000",
		16#02b5# => X"00000000",
		16#02b6# => X"00000000",
		16#02b7# => X"00000000",
		16#02b8# => X"00000000",
		16#02b9# => X"00000000",
		16#02ba# => X"00000000",
		16#02bb# => X"00000000",
		16#02bc# => X"00000000",
		16#02bd# => X"00000000",
		16#02be# => X"00000000",
		16#02bf# => X"00000000",
		16#02c0# => X"00000000",
		16#02c1# => X"00000000",
		16#02c2# => X"00000000",
		16#02c3# => X"00000000",
		16#02c4# => X"00000000",
		16#02c5# => X"00000000",
		16#02c6# => X"00000000",
		16#02c7# => X"00000000",
		16#02c8# => X"00000000",
		16#02c9# => X"00000000",
		16#02ca# => X"00000000",
		16#02cb# => X"00000000",
		16#02cc# => X"00000000",
		16#02cd# => X"00000000",
		16#02ce# => X"00000000",
		16#02cf# => X"00000000",
		16#02d0# => X"00000000",
		16#02d1# => X"00000000",
		16#02d2# => X"00000000",
		16#02d3# => X"00000000",
		16#02d4# => X"00000000",
		16#02d5# => X"00000000",
		16#02d6# => X"00000000",
		16#02d7# => X"00000000",
		16#02d8# => X"00000000",
		16#02d9# => X"00000000",
		16#02da# => X"00000000",
		16#02db# => X"00000000",
		16#02dc# => X"00000000",
		16#02dd# => X"00000000",
		16#02de# => X"00000000",
		16#02df# => X"00000000",
		16#02e0# => X"00000000",
		16#02e1# => X"00000000",
		16#02e2# => X"00000000",
		16#02e3# => X"00000000",
		16#02e4# => X"00000000",
		16#02e5# => X"00000000",
		16#02e6# => X"00000000",
		16#02e7# => X"00000000",
		16#02e8# => X"00000000",
		16#02e9# => X"00000000",
		16#02ea# => X"00000000",
		16#02eb# => X"00000000",
		16#02ec# => X"00000000",
		16#02ed# => X"00000000",
		16#02ee# => X"00000000",
		16#02ef# => X"00000000",
		16#02f0# => X"00000000",
		16#02f1# => X"00000000",
		16#02f2# => X"00000000",
		16#02f3# => X"00000000",
		16#02f4# => X"00000000",
		16#02f5# => X"00000000",
		16#02f6# => X"00000000",
		16#02f7# => X"00000000",
		16#02f8# => X"00000000",
		16#02f9# => X"00000000",
		16#02fa# => X"00000000",
		16#02fb# => X"00000000",
		16#02fc# => X"00000000",
		16#02fd# => X"00000000",
		16#02fe# => X"00000000",
		16#02ff# => X"00000000",
		16#0300# => X"00000000",
		16#0301# => X"00000000",
		16#0302# => X"00000000",
		16#0303# => X"00000000",
		16#0304# => X"00000000",
		16#0305# => X"00000000",
		16#0306# => X"00000000",
		16#0307# => X"00000000",
		16#0308# => X"00000000",
		16#0309# => X"00000000",
		16#030a# => X"00000000",
		16#030b# => X"00000000",
		16#030c# => X"00000000",
		16#030d# => X"00000000",
		16#030e# => X"00000000",
		16#030f# => X"00000000",
		16#0310# => X"00000000",
		16#0311# => X"00000000",
		16#0312# => X"00000000",
		16#0313# => X"00000000",
		16#0314# => X"00000000",
		16#0315# => X"00000000",
		16#0316# => X"00000000",
		16#0317# => X"00000000",
		16#0318# => X"00000000",
		16#0319# => X"00000000",
		16#031a# => X"00000000",
		16#031b# => X"00000000",
		16#031c# => X"00000000",
		16#031d# => X"00000000",
		16#031e# => X"00000000",
		16#031f# => X"00000000",
		16#0320# => X"00000000",
		16#0321# => X"00000000",
		16#0322# => X"00000000",
		16#0323# => X"00000000",
		16#0324# => X"00000000",
		16#0325# => X"00000000",
		16#0326# => X"00000000",
		16#0327# => X"00000000",
		16#0328# => X"00000000",
		16#0329# => X"00000000",
		16#032a# => X"00000000",
		16#032b# => X"00000000",
		16#032c# => X"00000000",
		16#032d# => X"00000000",
		16#032e# => X"00000000",
		16#032f# => X"00000000",
		16#0330# => X"00000000",
		16#0331# => X"00000000",
		16#0332# => X"00000000",
		16#0333# => X"00000000",
		16#0334# => X"00000000",
		16#0335# => X"00000000",
		16#0336# => X"00000000",
		16#0337# => X"00000000",
		16#0338# => X"00000000",
		16#0339# => X"00000000",
		16#033a# => X"00000000",
		16#033b# => X"00000000",
		16#033c# => X"00000000",
		16#033d# => X"00000000",
		16#033e# => X"00000000",
		16#033f# => X"00000000",
		16#0340# => X"00000000",
		16#0341# => X"00000000",
		16#0342# => X"00000000",
		16#0343# => X"00000000",
		16#0344# => X"00000000",
		16#0345# => X"00000000",
		16#0346# => X"00000000",
		16#0347# => X"00000000",
		16#0348# => X"00000000",
		16#0349# => X"00000000",
		16#034a# => X"00000000",
		16#034b# => X"00000000",
		16#034c# => X"00000000",
		16#034d# => X"00000000",
		16#034e# => X"00000000",
		16#034f# => X"00000000",
		16#0350# => X"00000000",
		16#0351# => X"00000000",
		16#0352# => X"00000000",
		16#0353# => X"00000000",
		16#0354# => X"00000000",
		16#0355# => X"00000000",
		16#0356# => X"00000000",
		16#0357# => X"00000000",
		16#0358# => X"00000000",
		16#0359# => X"00000000",
		16#035a# => X"00000000",
		16#035b# => X"00000000",
		16#035c# => X"00000000",
		16#035d# => X"00000000",
		16#035e# => X"00000000",
		16#035f# => X"00000000",
		16#0360# => X"00000000",
		16#0361# => X"00000000",
		16#0362# => X"00000000",
		16#0363# => X"00000000",
		16#0364# => X"00000000",
		16#0365# => X"00000000",
		16#0366# => X"00000000",
		16#0367# => X"00000000",
		16#0368# => X"00000000",
		16#0369# => X"00000000",
		16#036a# => X"00000000",
		16#036b# => X"00000000",
		16#036c# => X"00000000",
		16#036d# => X"00000000",
		16#036e# => X"00000000",
		16#036f# => X"00000000",
		16#0370# => X"00000000",
		16#0371# => X"00000000",
		16#0372# => X"00000000",
		16#0373# => X"00000000",
		16#0374# => X"00000000",
		16#0375# => X"00000000",
		16#0376# => X"00000000",
		16#0377# => X"00000000",
		16#0378# => X"00000000",
		16#0379# => X"00000000",
		16#037a# => X"00000000",
		16#037b# => X"00000000",
		16#037c# => X"00000000",
		16#037d# => X"00000000",
		16#037e# => X"00000000",
		16#037f# => X"00000000",
		16#0380# => X"00000000",
		16#0381# => X"00000000",
		16#0382# => X"00000000",
		16#0383# => X"00000000",
		16#0384# => X"00000000",
		16#0385# => X"00000000",
		16#0386# => X"00000000",
		16#0387# => X"00000000",
		16#0388# => X"00000000",
		16#0389# => X"00000000",
		16#038a# => X"00000000",
		16#038b# => X"00000000",
		16#038c# => X"00000000",
		16#038d# => X"00000000",
		16#038e# => X"00000000",
		16#038f# => X"00000000",
		16#0390# => X"00000000",
		16#0391# => X"00000000",
		16#0392# => X"00000000",
		16#0393# => X"00000000",
		16#0394# => X"00000000",
		16#0395# => X"00000000",
		16#0396# => X"00000000",
		16#0397# => X"00000000",
		16#0398# => X"00000000",
		16#0399# => X"00000000",
		16#039a# => X"00000000",
		16#039b# => X"00000000",
		16#039c# => X"00000000",
		16#039d# => X"00000000",
		16#039e# => X"00000000",
		16#039f# => X"00000000",
		16#03a0# => X"00000000",
		16#03a1# => X"00000000",
		16#03a2# => X"00000000",
		16#03a3# => X"00000000",
		16#03a4# => X"00000000",
		16#03a5# => X"00000000",
		16#03a6# => X"00000000",
		16#03a7# => X"00000000",
		16#03a8# => X"00000000",
		16#03a9# => X"00000000",
		16#03aa# => X"00000000",
		16#03ab# => X"00000000",
		16#03ac# => X"00000000",
		16#03ad# => X"00000000",
		16#03ae# => X"00000000",
		16#03af# => X"00000000",
		16#03b0# => X"00000000",
		16#03b1# => X"00000000",
		16#03b2# => X"00000000",
		16#03b3# => X"00000000",
		16#03b4# => X"00000000",
		16#03b5# => X"00000000",
		16#03b6# => X"00000000",
		16#03b7# => X"00000000",
		16#03b8# => X"00000000",
		16#03b9# => X"00000000",
		16#03ba# => X"00000000",
		16#03bb# => X"00000000",
		16#03bc# => X"00000000",
		16#03bd# => X"00000000",
		16#03be# => X"00000000",
		16#03bf# => X"00000000",
		16#03c0# => X"00000000",
		16#03c1# => X"00000000",
		16#03c2# => X"00000000",
		16#03c3# => X"00000000",
		16#03c4# => X"00000000",
		16#03c5# => X"00000000",
		16#03c6# => X"00000000",
		16#03c7# => X"00000000",
		16#03c8# => X"00000000",
		16#03c9# => X"00000000",
		16#03ca# => X"00000000",
		16#03cb# => X"00000000",
		16#03cc# => X"00000000",
		16#03cd# => X"00000000",
		16#03ce# => X"00000000",
		16#03cf# => X"00000000",
		16#03d0# => X"00000000",
		16#03d1# => X"00000000",
		16#03d2# => X"00000000",
		16#03d3# => X"00000000",
		16#03d4# => X"00000000",
		16#03d5# => X"00000000",
		16#03d6# => X"00000000",
		16#03d7# => X"00000000",
		16#03d8# => X"00000000",
		16#03d9# => X"00000000",
		16#03da# => X"00000000",
		16#03db# => X"00000000",
		16#03dc# => X"00000000",
		16#03dd# => X"00000000",
		16#03de# => X"00000000",
		16#03df# => X"00000000",
		16#03e0# => X"00000000",
		16#03e1# => X"00000000",
		16#03e2# => X"00000000",
		16#03e3# => X"00000000",
		16#03e4# => X"00000000",
		16#03e5# => X"00000000",
		16#03e6# => X"00000000",
		16#03e7# => X"00000000",
		16#03e8# => X"00000000",
		16#03e9# => X"00000000",
		16#03ea# => X"00000000",
		16#03eb# => X"00000000",
		16#03ec# => X"00000000",
		16#03ed# => X"00000000",
		16#03ee# => X"00000000",
		16#03ef# => X"00000000",
		16#03f0# => X"00000000",
		16#03f1# => X"00000000",
		16#03f2# => X"00000000",
		16#03f3# => X"00000000",
		16#03f4# => X"00000000",
		16#03f5# => X"00000000",
		16#03f6# => X"00000000",
		16#03f7# => X"00000000",
		16#03f8# => X"00000000",
		16#03f9# => X"00000000",
		16#03fa# => X"00000000",
		16#03fb# => X"00000000",
		16#03fc# => X"00000000",
		16#03fd# => X"00000000",
		16#03fe# => X"00000000",
		16#03ff# => X"00000000",
		16#0400# => X"f32e2034",
		16#0401# => X"13ce0e00",
		16#0402# => X"6302c003",
		16#0403# => X"13ce2e00",
		16#0404# => X"6300c005",
		16#0405# => X"13ce4e00",
		16#0406# => X"630ec005",
		16#0407# => X"13ce6e00",
		16#0408# => X"630cc007",
		16#0409# => X"13ce0e01",
		16#040a# => X"630ac009",
		16#040b# => X"971e0000",
		16#040c# => X"938e0e01",
		16#040d# => X"03ae0e00",
		16#040e# => X"130e1e00",
		16#040f# => X"23a0ce01",
		16#0410# => X"732e1034",
		16#0411# => X"130e4e00",
		16#0412# => X"73101e34",
		16#0413# => X"73002030",
		16#0414# => X"971e0000",
		16#0415# => X"938e0efe",
		16#0416# => X"03ae0e00",
		16#0417# => X"130e1e00",
		16#0418# => X"23a0ce01",
		16#0419# => X"732e1034",
		16#041a# => X"130e4e00",
		16#041b# => X"73101e34",
		16#041c# => X"73002030",
		16#041d# => X"971e0000",
		16#041e# => X"938e0efc",
		16#041f# => X"03ae0e00",
		16#0420# => X"130e1e00",
		16#0421# => X"23a0ce01",
		16#0422# => X"732e1034",
		16#0423# => X"130e4e00",
		16#0424# => X"73101e34",
		16#0425# => X"73002030",
		16#0426# => X"971e0000",
		16#0427# => X"938e0efa",
		16#0428# => X"03ae0e00",
		16#0429# => X"130e1e00",
		16#042a# => X"23a0ce01",
		16#042b# => X"732e1034",
		16#042c# => X"130e4e00",
		16#042d# => X"73101e34",
		16#042e# => X"73002030",
		16#042f# => X"971e0000",
		16#0430# => X"938e4ef8",
		16#0431# => X"03ae0e00",
		16#0432# => X"130e1e00",
		16#0433# => X"23a0ce01",
		16#0434# => X"f32e20fc",
		16#0435# => X"130e1000",
		16#0436# => X"93de1e00",
		16#0437# => X"93fc1e00",
		16#0438# => X"131e1e00",
		16#0439# => X"e38a0cfe",
		16#043a# => X"73200e7c",
		16#043b# => X"73002030",
		16#043c# => X"00000000",
		16#043d# => X"00000000",
		16#043e# => X"00000000",
		16#043f# => X"00000000",
		16#0440# => X"00000000",
		16#0441# => X"00000000",
		16#0442# => X"00000000",
		16#0443# => X"00000000",
		16#0444# => X"00000000",
		16#0445# => X"00000000",
		16#0446# => X"00000000",
		16#0447# => X"00000000",
		16#0448# => X"00000000",
		16#0449# => X"00000000",
		16#044a# => X"00000000",
		16#044b# => X"00000000",
		16#044c# => X"00000000",
		16#044d# => X"00000000",
		16#044e# => X"00000000",
		16#044f# => X"00000000",
		16#0450# => X"00000000",
		16#0451# => X"00000000",
		16#0452# => X"00000000",
		16#0453# => X"00000000",
		16#0454# => X"00000000",
		16#0455# => X"00000000",
		16#0456# => X"00000000",
		16#0457# => X"00000000",
		16#0458# => X"00000000",
		16#0459# => X"00000000",
		16#045a# => X"00000000",
		16#045b# => X"00000000",
		16#045c# => X"00000000",
		16#045d# => X"00000000",
		16#045e# => X"00000000",
		16#045f# => X"00000000",
		16#0460# => X"00000000",
		16#0461# => X"00000000",
		16#0462# => X"00000000",
		16#0463# => X"00000000",
		16#0464# => X"00000000",
		16#0465# => X"00000000",
		16#0466# => X"00000000",
		16#0467# => X"00000000",
		16#0468# => X"00000000",
		16#0469# => X"00000000",
		16#046a# => X"00000000",
		16#046b# => X"00000000",
		16#046c# => X"00000000",
		16#046d# => X"00000000",
		16#046e# => X"00000000",
		16#046f# => X"00000000",
		16#0470# => X"00000000",
		16#0471# => X"00000000",
		16#0472# => X"00000000",
		16#0473# => X"00000000",
		16#0474# => X"00000000",
		16#0475# => X"00000000",
		16#0476# => X"00000000",
		16#0477# => X"00000000",
		16#0478# => X"00000000",
		16#0479# => X"00000000",
		16#047a# => X"00000000",
		16#047b# => X"00000000",
		16#047c# => X"00000000",
		16#047d# => X"00000000",
		16#047e# => X"00000000",
		16#047f# => X"00000000",
		16#0480# => X"00000000",
		16#0481# => X"00000000",
		16#0482# => X"00000000",
		16#0483# => X"00000000",
		16#0484# => X"00000000",
		16#0485# => X"00000000",
		16#0486# => X"00000000",
		16#0487# => X"00000000",
		16#0488# => X"00000000",
		16#0489# => X"00000000",
		16#048a# => X"00000000",
		16#048b# => X"00000000",
		16#048c# => X"00000000",
		16#048d# => X"00000000",
		16#048e# => X"00000000",
		16#048f# => X"00000000",
		16#0490# => X"00000000",
		16#0491# => X"00000000",
		16#0492# => X"00000000",
		16#0493# => X"00000000",
		16#0494# => X"00000000",
		16#0495# => X"00000000",
		16#0496# => X"00000000",
		16#0497# => X"00000000",
		16#0498# => X"00000000",
		16#0499# => X"00000000",
		16#049a# => X"00000000",
		16#049b# => X"00000000",
		16#049c# => X"00000000",
		16#049d# => X"00000000",
		16#049e# => X"00000000",
		16#049f# => X"00000000",
		16#04a0# => X"00000000",
		16#04a1# => X"00000000",
		16#04a2# => X"00000000",
		16#04a3# => X"00000000",
		16#04a4# => X"00000000",
		16#04a5# => X"00000000",
		16#04a6# => X"00000000",
		16#04a7# => X"00000000",
		16#04a8# => X"00000000",
		16#04a9# => X"00000000",
		16#04aa# => X"00000000",
		16#04ab# => X"00000000",
		16#04ac# => X"00000000",
		16#04ad# => X"00000000",
		16#04ae# => X"00000000",
		16#04af# => X"00000000",
		16#04b0# => X"00000000",
		16#04b1# => X"00000000",
		16#04b2# => X"00000000",
		16#04b3# => X"00000000",
		16#04b4# => X"00000000",
		16#04b5# => X"00000000",
		16#04b6# => X"00000000",
		16#04b7# => X"00000000",
		16#04b8# => X"00000000",
		16#04b9# => X"00000000",
		16#04ba# => X"00000000",
		16#04bb# => X"00000000",
		16#04bc# => X"00000000",
		16#04bd# => X"00000000",
		16#04be# => X"00000000",
		16#04bf# => X"00000000",
		16#04c0# => X"00000000",
		16#04c1# => X"00000000",
		16#04c2# => X"00000000",
		16#04c3# => X"00000000",
		16#04c4# => X"00000000",
		16#04c5# => X"00000000",
		16#04c6# => X"00000000",
		16#04c7# => X"00000000",
		16#04c8# => X"00000000",
		16#04c9# => X"00000000",
		16#04ca# => X"00000000",
		16#04cb# => X"00000000",
		16#04cc# => X"00000000",
		16#04cd# => X"00000000",
		16#04ce# => X"00000000",
		16#04cf# => X"00000000",
		16#04d0# => X"00000000",
		16#04d1# => X"00000000",
		16#04d2# => X"00000000",
		16#04d3# => X"00000000",
		16#04d4# => X"00000000",
		16#04d5# => X"00000000",
		16#04d6# => X"00000000",
		16#04d7# => X"00000000",
		16#04d8# => X"00000000",
		16#04d9# => X"00000000",
		16#04da# => X"00000000",
		16#04db# => X"00000000",
		16#04dc# => X"00000000",
		16#04dd# => X"00000000",
		16#04de# => X"00000000",
		16#04df# => X"00000000",
		16#04e0# => X"00000000",
		16#04e1# => X"00000000",
		16#04e2# => X"00000000",
		16#04e3# => X"00000000",
		16#04e4# => X"00000000",
		16#04e5# => X"00000000",
		16#04e6# => X"00000000",
		16#04e7# => X"00000000",
		16#04e8# => X"00000000",
		16#04e9# => X"00000000",
		16#04ea# => X"00000000",
		16#04eb# => X"00000000",
		16#04ec# => X"00000000",
		16#04ed# => X"00000000",
		16#04ee# => X"00000000",
		16#04ef# => X"00000000",
		16#04f0# => X"00000000",
		16#04f1# => X"00000000",
		16#04f2# => X"00000000",
		16#04f3# => X"00000000",
		16#04f4# => X"00000000",
		16#04f5# => X"00000000",
		16#04f6# => X"00000000",
		16#04f7# => X"00000000",
		16#04f8# => X"00000000",
		16#04f9# => X"00000000",
		16#04fa# => X"00000000",
		16#04fb# => X"00000000",
		16#04fc# => X"00000000",
		16#04fd# => X"00000000",
		16#04fe# => X"00000000",
		16#04ff# => X"00000000",
		16#0500# => X"00000000",
		16#0501# => X"00000000",
		16#0502# => X"00000000",
		16#0503# => X"00000000",
		16#0504# => X"00000000",
		16#0505# => X"00000000",
		16#0506# => X"00000000",
		16#0507# => X"00000000",
		16#0508# => X"00000000",
		16#0509# => X"00000000",
		16#050a# => X"00000000",
		16#050b# => X"00000000",
		16#050c# => X"00000000",
		16#050d# => X"00000000",
		16#050e# => X"00000000",
		16#050f# => X"00000000",
		16#0510# => X"00000000",
		16#0511# => X"00000000",
		16#0512# => X"00000000",
		16#0513# => X"00000000",
		16#0514# => X"00000000",
		16#0515# => X"00000000",
		16#0516# => X"00000000",
		16#0517# => X"00000000",
		16#0518# => X"00000000",
		16#0519# => X"00000000",
		16#051a# => X"00000000",
		16#051b# => X"00000000",
		16#051c# => X"00000000",
		16#051d# => X"00000000",
		16#051e# => X"00000000",
		16#051f# => X"00000000",
		16#0520# => X"00000000",
		16#0521# => X"00000000",
		16#0522# => X"00000000",
		16#0523# => X"00000000",
		16#0524# => X"00000000",
		16#0525# => X"00000000",
		16#0526# => X"00000000",
		16#0527# => X"00000000",
		16#0528# => X"00000000",
		16#0529# => X"00000000",
		16#052a# => X"00000000",
		16#052b# => X"00000000",
		16#052c# => X"00000000",
		16#052d# => X"00000000",
		16#052e# => X"00000000",
		16#052f# => X"00000000",
		16#0530# => X"00000000",
		16#0531# => X"00000000",
		16#0532# => X"00000000",
		16#0533# => X"00000000",
		16#0534# => X"00000000",
		16#0535# => X"00000000",
		16#0536# => X"00000000",
		16#0537# => X"00000000",
		16#0538# => X"00000000",
		16#0539# => X"00000000",
		16#053a# => X"00000000",
		16#053b# => X"00000000",
		16#053c# => X"00000000",
		16#053d# => X"00000000",
		16#053e# => X"00000000",
		16#053f# => X"00000000",
		16#0540# => X"00000000",
		16#0541# => X"00000000",
		16#0542# => X"00000000",
		16#0543# => X"00000000",
		16#0544# => X"00000000",
		16#0545# => X"00000000",
		16#0546# => X"00000000",
		16#0547# => X"00000000",
		16#0548# => X"00000000",
		16#0549# => X"00000000",
		16#054a# => X"00000000",
		16#054b# => X"00000000",
		16#054c# => X"00000000",
		16#054d# => X"00000000",
		16#054e# => X"00000000",
		16#054f# => X"00000000",
		16#0550# => X"00000000",
		16#0551# => X"00000000",
		16#0552# => X"00000000",
		16#0553# => X"00000000",
		16#0554# => X"00000000",
		16#0555# => X"00000000",
		16#0556# => X"00000000",
		16#0557# => X"00000000",
		16#0558# => X"00000000",
		16#0559# => X"00000000",
		16#055a# => X"00000000",
		16#055b# => X"00000000",
		16#055c# => X"00000000",
		16#055d# => X"00000000",
		16#055e# => X"00000000",
		16#055f# => X"00000000",
		16#0560# => X"00000000",
		16#0561# => X"00000000",
		16#0562# => X"00000000",
		16#0563# => X"00000000",
		16#0564# => X"00000000",
		16#0565# => X"00000000",
		16#0566# => X"00000000",
		16#0567# => X"00000000",
		16#0568# => X"00000000",
		16#0569# => X"00000000",
		16#056a# => X"00000000",
		16#056b# => X"00000000",
		16#056c# => X"00000000",
		16#056d# => X"00000000",
		16#056e# => X"00000000",
		16#056f# => X"00000000",
		16#0570# => X"00000000",
		16#0571# => X"00000000",
		16#0572# => X"00000000",
		16#0573# => X"00000000",
		16#0574# => X"00000000",
		16#0575# => X"00000000",
		16#0576# => X"00000000",
		16#0577# => X"00000000",
		16#0578# => X"00000000",
		16#0579# => X"00000000",
		16#057a# => X"00000000",
		16#057b# => X"00000000",
		16#057c# => X"00000000",
		16#057d# => X"00000000",
		16#057e# => X"00000000",
		16#057f# => X"00000000",
		16#0580# => X"00000000",
		16#0581# => X"00000000",
		16#0582# => X"00000000",
		16#0583# => X"00000000",
		16#0584# => X"00000000",
		16#0585# => X"00000000",
		16#0586# => X"00000000",
		16#0587# => X"00000000",
		16#0588# => X"00000000",
		16#0589# => X"00000000",
		16#058a# => X"00000000",
		16#058b# => X"00000000",
		16#058c# => X"00000000",
		16#058d# => X"00000000",
		16#058e# => X"00000000",
		16#058f# => X"00000000",
		16#0590# => X"00000000",
		16#0591# => X"00000000",
		16#0592# => X"00000000",
		16#0593# => X"00000000",
		16#0594# => X"00000000",
		16#0595# => X"00000000",
		16#0596# => X"00000000",
		16#0597# => X"00000000",
		16#0598# => X"00000000",
		16#0599# => X"00000000",
		16#059a# => X"00000000",
		16#059b# => X"00000000",
		16#059c# => X"00000000",
		16#059d# => X"00000000",
		16#059e# => X"00000000",
		16#059f# => X"00000000",
		16#05a0# => X"00000000",
		16#05a1# => X"00000000",
		16#05a2# => X"00000000",
		16#05a3# => X"00000000",
		16#05a4# => X"00000000",
		16#05a5# => X"00000000",
		16#05a6# => X"00000000",
		16#05a7# => X"00000000",
		16#05a8# => X"00000000",
		16#05a9# => X"00000000",
		16#05aa# => X"00000000",
		16#05ab# => X"00000000",
		16#05ac# => X"00000000",
		16#05ad# => X"00000000",
		16#05ae# => X"00000000",
		16#05af# => X"00000000",
		16#05b0# => X"00000000",
		16#05b1# => X"00000000",
		16#05b2# => X"00000000",
		16#05b3# => X"00000000",
		16#05b4# => X"00000000",
		16#05b5# => X"00000000",
		16#05b6# => X"00000000",
		16#05b7# => X"00000000",
		16#05b8# => X"00000000",
		16#05b9# => X"00000000",
		16#05ba# => X"00000000",
		16#05bb# => X"00000000",
		16#05bc# => X"00000000",
		16#05bd# => X"00000000",
		16#05be# => X"00000000",
		16#05bf# => X"00000000",
		16#05c0# => X"00000000",
		16#05c1# => X"00000000",
		16#05c2# => X"00000000",
		16#05c3# => X"00000000",
		16#05c4# => X"00000000",
		16#05c5# => X"00000000",
		16#05c6# => X"00000000",
		16#05c7# => X"00000000",
		16#05c8# => X"00000000",
		16#05c9# => X"00000000",
		16#05ca# => X"00000000",
		16#05cb# => X"00000000",
		16#05cc# => X"00000000",
		16#05cd# => X"00000000",
		16#05ce# => X"00000000",
		16#05cf# => X"00000000",
		16#05d0# => X"00000000",
		16#05d1# => X"00000000",
		16#05d2# => X"00000000",
		16#05d3# => X"00000000",
		16#05d4# => X"00000000",
		16#05d5# => X"00000000",
		16#05d6# => X"00000000",
		16#05d7# => X"00000000",
		16#05d8# => X"00000000",
		16#05d9# => X"00000000",
		16#05da# => X"00000000",
		16#05db# => X"00000000",
		16#05dc# => X"00000000",
		16#05dd# => X"00000000",
		16#05de# => X"00000000",
		16#05df# => X"00000000",
		16#05e0# => X"00000000",
		16#05e1# => X"00000000",
		16#05e2# => X"00000000",
		16#05e3# => X"00000000",
		16#05e4# => X"00000000",
		16#05e5# => X"00000000",
		16#05e6# => X"00000000",
		16#05e7# => X"00000000",
		16#05e8# => X"00000000",
		16#05e9# => X"00000000",
		16#05ea# => X"00000000",
		16#05eb# => X"00000000",
		16#05ec# => X"00000000",
		16#05ed# => X"00000000",
		16#05ee# => X"00000000",
		16#05ef# => X"00000000",
		16#05f0# => X"00000000",
		16#05f1# => X"00000000",
		16#05f2# => X"00000000",
		16#05f3# => X"00000000",
		16#05f4# => X"00000000",
		16#05f5# => X"00000000",
		16#05f6# => X"00000000",
		16#05f7# => X"00000000",
		16#05f8# => X"00000000",
		16#05f9# => X"00000000",
		16#05fa# => X"00000000",
		16#05fb# => X"00000000",
		16#05fc# => X"00000000",
		16#05fd# => X"00000000",
		16#05fe# => X"00000000",
		16#05ff# => X"00000000",
		16#0600# => X"00000000",
		16#0601# => X"00000000",
		16#0602# => X"00000000",
		16#0603# => X"00000000",
		16#0604# => X"00000000",
		16#0605# => X"00000000",
		16#0606# => X"00000000",
		16#0607# => X"00000000",
		16#0608# => X"00000000",
		16#0609# => X"00000000",
		16#060a# => X"00000000",
		16#060b# => X"00000000",
		16#060c# => X"00000000",
		16#060d# => X"00000000",
		16#060e# => X"00000000",
		16#060f# => X"00000000",
		16#0610# => X"00000000",
		16#0611# => X"00000000",
		16#0612# => X"00000000",
		16#0613# => X"00000000",
		16#0614# => X"00000000",
		16#0615# => X"00000000",
		16#0616# => X"00000000",
		16#0617# => X"00000000",
		16#0618# => X"00000000",
		16#0619# => X"00000000",
		16#061a# => X"00000000",
		16#061b# => X"00000000",
		16#061c# => X"00000000",
		16#061d# => X"00000000",
		16#061e# => X"00000000",
		16#061f# => X"00000000",
		16#0620# => X"00000000",
		16#0621# => X"00000000",
		16#0622# => X"00000000",
		16#0623# => X"00000000",
		16#0624# => X"00000000",
		16#0625# => X"00000000",
		16#0626# => X"00000000",
		16#0627# => X"00000000",
		16#0628# => X"00000000",
		16#0629# => X"00000000",
		16#062a# => X"00000000",
		16#062b# => X"00000000",
		16#062c# => X"00000000",
		16#062d# => X"00000000",
		16#062e# => X"00000000",
		16#062f# => X"00000000",
		16#0630# => X"00000000",
		16#0631# => X"00000000",
		16#0632# => X"00000000",
		16#0633# => X"00000000",
		16#0634# => X"00000000",
		16#0635# => X"00000000",
		16#0636# => X"00000000",
		16#0637# => X"00000000",
		16#0638# => X"00000000",
		16#0639# => X"00000000",
		16#063a# => X"00000000",
		16#063b# => X"00000000",
		16#063c# => X"00000000",
		16#063d# => X"00000000",
		16#063e# => X"00000000",
		16#063f# => X"00000000",
		16#0640# => X"00000000",
		16#0641# => X"00000000",
		16#0642# => X"00000000",
		16#0643# => X"00000000",
		16#0644# => X"00000000",
		16#0645# => X"00000000",
		16#0646# => X"00000000",
		16#0647# => X"00000000",
		16#0648# => X"00000000",
		16#0649# => X"00000000",
		16#064a# => X"00000000",
		16#064b# => X"00000000",
		16#064c# => X"00000000",
		16#064d# => X"00000000",
		16#064e# => X"00000000",
		16#064f# => X"00000000",
		16#0650# => X"00000000",
		16#0651# => X"00000000",
		16#0652# => X"00000000",
		16#0653# => X"00000000",
		16#0654# => X"00000000",
		16#0655# => X"00000000",
		16#0656# => X"00000000",
		16#0657# => X"00000000",
		16#0658# => X"00000000",
		16#0659# => X"00000000",
		16#065a# => X"00000000",
		16#065b# => X"00000000",
		16#065c# => X"00000000",
		16#065d# => X"00000000",
		16#065e# => X"00000000",
		16#065f# => X"00000000",
		16#0660# => X"00000000",
		16#0661# => X"00000000",
		16#0662# => X"00000000",
		16#0663# => X"00000000",
		16#0664# => X"00000000",
		16#0665# => X"00000000",
		16#0666# => X"00000000",
		16#0667# => X"00000000",
		16#0668# => X"00000000",
		16#0669# => X"00000000",
		16#066a# => X"00000000",
		16#066b# => X"00000000",
		16#066c# => X"00000000",
		16#066d# => X"00000000",
		16#066e# => X"00000000",
		16#066f# => X"00000000",
		16#0670# => X"00000000",
		16#0671# => X"00000000",
		16#0672# => X"00000000",
		16#0673# => X"00000000",
		16#0674# => X"00000000",
		16#0675# => X"00000000",
		16#0676# => X"00000000",
		16#0677# => X"00000000",
		16#0678# => X"00000000",
		16#0679# => X"00000000",
		16#067a# => X"00000000",
		16#067b# => X"00000000",
		16#067c# => X"00000000",
		16#067d# => X"00000000",
		16#067e# => X"00000000",
		16#067f# => X"00000000",
		16#0680# => X"00000000",
		16#0681# => X"00000000",
		16#0682# => X"00000000",
		16#0683# => X"00000000",
		16#0684# => X"00000000",
		16#0685# => X"00000000",
		16#0686# => X"00000000",
		16#0687# => X"00000000",
		16#0688# => X"00000000",
		16#0689# => X"00000000",
		16#068a# => X"00000000",
		16#068b# => X"00000000",
		16#068c# => X"00000000",
		16#068d# => X"00000000",
		16#068e# => X"00000000",
		16#068f# => X"00000000",
		16#0690# => X"00000000",
		16#0691# => X"00000000",
		16#0692# => X"00000000",
		16#0693# => X"00000000",
		16#0694# => X"00000000",
		16#0695# => X"00000000",
		16#0696# => X"00000000",
		16#0697# => X"00000000",
		16#0698# => X"00000000",
		16#0699# => X"00000000",
		16#069a# => X"00000000",
		16#069b# => X"00000000",
		16#069c# => X"00000000",
		16#069d# => X"00000000",
		16#069e# => X"00000000",
		16#069f# => X"00000000",
		16#06a0# => X"00000000",
		16#06a1# => X"00000000",
		16#06a2# => X"00000000",
		16#06a3# => X"00000000",
		16#06a4# => X"00000000",
		16#06a5# => X"00000000",
		16#06a6# => X"00000000",
		16#06a7# => X"00000000",
		16#06a8# => X"00000000",
		16#06a9# => X"00000000",
		16#06aa# => X"00000000",
		16#06ab# => X"00000000",
		16#06ac# => X"00000000",
		16#06ad# => X"00000000",
		16#06ae# => X"00000000",
		16#06af# => X"00000000",
		16#06b0# => X"00000000",
		16#06b1# => X"00000000",
		16#06b2# => X"00000000",
		16#06b3# => X"00000000",
		16#06b4# => X"00000000",
		16#06b5# => X"00000000",
		16#06b6# => X"00000000",
		16#06b7# => X"00000000",
		16#06b8# => X"00000000",
		16#06b9# => X"00000000",
		16#06ba# => X"00000000",
		16#06bb# => X"00000000",
		16#06bc# => X"00000000",
		16#06bd# => X"00000000",
		16#06be# => X"00000000",
		16#06bf# => X"00000000",
		16#06c0# => X"00000000",
		16#06c1# => X"00000000",
		16#06c2# => X"00000000",
		16#06c3# => X"00000000",
		16#06c4# => X"00000000",
		16#06c5# => X"00000000",
		16#06c6# => X"00000000",
		16#06c7# => X"00000000",
		16#06c8# => X"00000000",
		16#06c9# => X"00000000",
		16#06ca# => X"00000000",
		16#06cb# => X"00000000",
		16#06cc# => X"00000000",
		16#06cd# => X"00000000",
		16#06ce# => X"00000000",
		16#06cf# => X"00000000",
		16#06d0# => X"00000000",
		16#06d1# => X"00000000",
		16#06d2# => X"00000000",
		16#06d3# => X"00000000",
		16#06d4# => X"00000000",
		16#06d5# => X"00000000",
		16#06d6# => X"00000000",
		16#06d7# => X"00000000",
		16#06d8# => X"00000000",
		16#06d9# => X"00000000",
		16#06da# => X"00000000",
		16#06db# => X"00000000",
		16#06dc# => X"00000000",
		16#06dd# => X"00000000",
		16#06de# => X"00000000",
		16#06df# => X"00000000",
		16#06e0# => X"00000000",
		16#06e1# => X"00000000",
		16#06e2# => X"00000000",
		16#06e3# => X"00000000",
		16#06e4# => X"00000000",
		16#06e5# => X"00000000",
		16#06e6# => X"00000000",
		16#06e7# => X"00000000",
		16#06e8# => X"00000000",
		16#06e9# => X"00000000",
		16#06ea# => X"00000000",
		16#06eb# => X"00000000",
		16#06ec# => X"00000000",
		16#06ed# => X"00000000",
		16#06ee# => X"00000000",
		16#06ef# => X"00000000",
		16#06f0# => X"00000000",
		16#06f1# => X"00000000",
		16#06f2# => X"00000000",
		16#06f3# => X"00000000",
		16#06f4# => X"00000000",
		16#06f5# => X"00000000",
		16#06f6# => X"00000000",
		16#06f7# => X"00000000",
		16#06f8# => X"00000000",
		16#06f9# => X"00000000",
		16#06fa# => X"00000000",
		16#06fb# => X"00000000",
		16#06fc# => X"00000000",
		16#06fd# => X"00000000",
		16#06fe# => X"00000000",
		16#06ff# => X"00000000",
		16#0700# => X"00000000",
		16#0701# => X"00000000",
		16#0702# => X"00000000",
		16#0703# => X"00000000",
		16#0704# => X"00000000",
		16#0705# => X"00000000",
		16#0706# => X"00000000",
		16#0707# => X"00000000",
		16#0708# => X"00000000",
		16#0709# => X"00000000",
		16#070a# => X"00000000",
		16#070b# => X"00000000",
		16#070c# => X"00000000",
		16#070d# => X"00000000",
		16#070e# => X"00000000",
		16#070f# => X"00000000",
		16#0710# => X"00000000",
		16#0711# => X"00000000",
		16#0712# => X"00000000",
		16#0713# => X"00000000",
		16#0714# => X"00000000",
		16#0715# => X"00000000",
		16#0716# => X"00000000",
		16#0717# => X"00000000",
		16#0718# => X"00000000",
		16#0719# => X"00000000",
		16#071a# => X"00000000",
		16#071b# => X"00000000",
		16#071c# => X"00000000",
		16#071d# => X"00000000",
		16#071e# => X"00000000",
		16#071f# => X"00000000",
		16#0720# => X"00000000",
		16#0721# => X"00000000",
		16#0722# => X"00000000",
		16#0723# => X"00000000",
		16#0724# => X"00000000",
		16#0725# => X"00000000",
		16#0726# => X"00000000",
		16#0727# => X"00000000",
		16#0728# => X"00000000",
		16#0729# => X"00000000",
		16#072a# => X"00000000",
		16#072b# => X"00000000",
		16#072c# => X"00000000",
		16#072d# => X"00000000",
		16#072e# => X"00000000",
		16#072f# => X"00000000",
		16#0730# => X"00000000",
		16#0731# => X"00000000",
		16#0732# => X"00000000",
		16#0733# => X"00000000",
		16#0734# => X"00000000",
		16#0735# => X"00000000",
		16#0736# => X"00000000",
		16#0737# => X"00000000",
		16#0738# => X"00000000",
		16#0739# => X"00000000",
		16#073a# => X"00000000",
		16#073b# => X"00000000",
		16#073c# => X"00000000",
		16#073d# => X"00000000",
		16#073e# => X"00000000",
		16#073f# => X"00000000",
		16#0740# => X"00000000",
		16#0741# => X"00000000",
		16#0742# => X"00000000",
		16#0743# => X"00000000",
		16#0744# => X"00000000",
		16#0745# => X"00000000",
		16#0746# => X"00000000",
		16#0747# => X"00000000",
		16#0748# => X"00000000",
		16#0749# => X"00000000",
		16#074a# => X"00000000",
		16#074b# => X"00000000",
		16#074c# => X"00000000",
		16#074d# => X"00000000",
		16#074e# => X"00000000",
		16#074f# => X"00000000",
		16#0750# => X"00000000",
		16#0751# => X"00000000",
		16#0752# => X"00000000",
		16#0753# => X"00000000",
		16#0754# => X"00000000",
		16#0755# => X"00000000",
		16#0756# => X"00000000",
		16#0757# => X"00000000",
		16#0758# => X"00000000",
		16#0759# => X"00000000",
		16#075a# => X"00000000",
		16#075b# => X"00000000",
		16#075c# => X"00000000",
		16#075d# => X"00000000",
		16#075e# => X"00000000",
		16#075f# => X"00000000",
		16#0760# => X"00000000",
		16#0761# => X"00000000",
		16#0762# => X"00000000",
		16#0763# => X"00000000",
		16#0764# => X"00000000",
		16#0765# => X"00000000",
		16#0766# => X"00000000",
		16#0767# => X"00000000",
		16#0768# => X"00000000",
		16#0769# => X"00000000",
		16#076a# => X"00000000",
		16#076b# => X"00000000",
		16#076c# => X"00000000",
		16#076d# => X"00000000",
		16#076e# => X"00000000",
		16#076f# => X"00000000",
		16#0770# => X"00000000",
		16#0771# => X"00000000",
		16#0772# => X"00000000",
		16#0773# => X"00000000",
		16#0774# => X"00000000",
		16#0775# => X"00000000",
		16#0776# => X"00000000",
		16#0777# => X"00000000",
		16#0778# => X"00000000",
		16#0779# => X"00000000",
		16#077a# => X"00000000",
		16#077b# => X"00000000",
		16#077c# => X"00000000",
		16#077d# => X"00000000",
		16#077e# => X"00000000",
		16#077f# => X"00000000",
		16#0780# => X"00000000",
		16#0781# => X"00000000",
		16#0782# => X"00000000",
		16#0783# => X"00000000",
		16#0784# => X"00000000",
		16#0785# => X"00000000",
		16#0786# => X"00000000",
		16#0787# => X"00000000",
		16#0788# => X"00000000",
		16#0789# => X"00000000",
		16#078a# => X"00000000",
		16#078b# => X"00000000",
		16#078c# => X"00000000",
		16#078d# => X"00000000",
		16#078e# => X"00000000",
		16#078f# => X"00000000",
		16#0790# => X"00000000",
		16#0791# => X"00000000",
		16#0792# => X"00000000",
		16#0793# => X"00000000",
		16#0794# => X"00000000",
		16#0795# => X"00000000",
		16#0796# => X"00000000",
		16#0797# => X"00000000",
		16#0798# => X"00000000",
		16#0799# => X"00000000",
		16#079a# => X"00000000",
		16#079b# => X"00000000",
		16#079c# => X"00000000",
		16#079d# => X"00000000",
		16#079e# => X"00000000",
		16#079f# => X"00000000",
		16#07a0# => X"00000000",
		16#07a1# => X"00000000",
		16#07a2# => X"00000000",
		16#07a3# => X"00000000",
		16#07a4# => X"00000000",
		16#07a5# => X"00000000",
		16#07a6# => X"00000000",
		16#07a7# => X"00000000",
		16#07a8# => X"00000000",
		16#07a9# => X"00000000",
		16#07aa# => X"00000000",
		16#07ab# => X"00000000",
		16#07ac# => X"00000000",
		16#07ad# => X"00000000",
		16#07ae# => X"00000000",
		16#07af# => X"00000000",
		16#07b0# => X"00000000",
		16#07b1# => X"00000000",
		16#07b2# => X"00000000",
		16#07b3# => X"00000000",
		16#07b4# => X"00000000",
		16#07b5# => X"00000000",
		16#07b6# => X"00000000",
		16#07b7# => X"00000000",
		16#07b8# => X"00000000",
		16#07b9# => X"00000000",
		16#07ba# => X"00000000",
		16#07bb# => X"00000000",
		16#07bc# => X"00000000",
		16#07bd# => X"00000000",
		16#07be# => X"00000000",
		16#07bf# => X"00000000",
		16#07c0# => X"00000000",
		16#07c1# => X"00000000",
		16#07c2# => X"00000000",
		16#07c3# => X"00000000",
		16#07c4# => X"00000000",
		16#07c5# => X"00000000",
		16#07c6# => X"00000000",
		16#07c7# => X"00000000",
		16#07c8# => X"00000000",
		16#07c9# => X"00000000",
		16#07ca# => X"00000000",
		16#07cb# => X"00000000",
		16#07cc# => X"00000000",
		16#07cd# => X"00000000",
		16#07ce# => X"00000000",
		16#07cf# => X"00000000",
		16#07d0# => X"00000000",
		16#07d1# => X"00000000",
		16#07d2# => X"00000000",
		16#07d3# => X"00000000",
		16#07d4# => X"00000000",
		16#07d5# => X"00000000",
		16#07d6# => X"00000000",
		16#07d7# => X"00000000",
		16#07d8# => X"00000000",
		16#07d9# => X"00000000",
		16#07da# => X"00000000",
		16#07db# => X"00000000",
		16#07dc# => X"00000000",
		16#07dd# => X"00000000",
		16#07de# => X"00000000",
		16#07df# => X"00000000",
		16#07e0# => X"00000000",
		16#07e1# => X"00000000",
		16#07e2# => X"00000000",
		16#07e3# => X"00000000",
		16#07e4# => X"00000000",
		16#07e5# => X"00000000",
		16#07e6# => X"00000000",
		16#07e7# => X"00000000",
		16#07e8# => X"00000000",
		16#07e9# => X"00000000",
		16#07ea# => X"00000000",
		16#07eb# => X"00000000",
		16#07ec# => X"00000000",
		16#07ed# => X"00000000",
		16#07ee# => X"00000000",
		16#07ef# => X"00000000",
		16#07f0# => X"00000000",
		16#07f1# => X"00000000",
		16#07f2# => X"00000000",
		16#07f3# => X"00000000",
		16#07f4# => X"00000000",
		16#07f5# => X"00000000",
		16#07f6# => X"00000000",
		16#07f7# => X"00000000",
		16#07f8# => X"00000000",
		16#07f9# => X"00000000",
		16#07fa# => X"00000000",
		16#07fb# => X"00000000",
		16#07fc# => X"00000000",
		16#07fd# => X"00000000",
		16#07fe# => X"00000000",
		16#07ff# => X"00000000",
		16#0800# => X"ffffffff",
		16#0801# => X"ffffffff",
		16#0802# => X"ffffffff",
		16#0803# => X"ffffffff",
		16#0804# => X"ffffffff",
		16#0805# => X"ffffffff",
		16#0806# => X"ffffffff",
		16#0807# => X"ffffffff",
		16#0808# => X"ffffffff",
		16#0809# => X"ffffffff",
		16#080a# => X"ffffffff",
		16#080b# => X"efbeadde",
		16#080c# => X"00000000",
		16#080d# => X"00000000",
		16#080e# => X"00000000",
		16#080f# => X"00000000",
		16#0810# => X"00000000",
		16#0811# => X"00000000",
		16#0812# => X"00000000",
		others => X"00000000"
	);

end package;